`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/23/2021 03:13:04 PM
// Design Name: 
// Module Name: DataMemory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module DataMemory(Address, WriteData, Clk, MemWrite, MemRead, ReadData, whb); 

    input [31:0] Address; 	                                 // Input Address 
    input [31:0] WriteData;                                  // Data that needs to be written into the address 
    input Clk;
    input MemWrite; 		                                 // Control signal for memory write 
    input MemRead; 			                                 // Control signal for memory read 
    input [1:0] whb;
    
    output reg[31:0] ReadData;                               // Contents of memory location at Address

    reg [31:0] memory [0:8191];
    
    initial begin
    //$readmemh("data_memory.mem",memory);
    
  memory[0] <= 32'h27;
memory[1] <= 32'h1f;
memory[2] <= 32'h8;
memory[3] <= 32'h4;
memory[4] <= 32'h0;
memory[5] <= 32'h0;
memory[6] <= 32'h0;
memory[7] <= 32'h0;
memory[8] <= 32'h0;
memory[9] <= 32'h0;
memory[10] <= 32'h0;
memory[11] <= 32'h0;
memory[12] <= 32'h0;
memory[13] <= 32'h0;
memory[14] <= 32'h0;
memory[15] <= 32'h0;
memory[16] <= 32'h0;
memory[17] <= 32'h0;
memory[18] <= 32'h0;
memory[19] <= 32'h0;
memory[20] <= 32'h0;
memory[21] <= 32'h0;
memory[22] <= 32'h0;
memory[23] <= 32'h0;
memory[24] <= 32'h0;
memory[25] <= 32'h0;
memory[26] <= 32'h0;
memory[27] <= 32'h0;
memory[28] <= 32'h0;
memory[29] <= 32'h0;
memory[30] <= 32'h0;
memory[31] <= 32'h1;
memory[32] <= 32'h1;
memory[33] <= 32'h1;
memory[34] <= 32'h1;
memory[35] <= 32'h0;
memory[36] <= 32'h0;
memory[37] <= 32'h0;
memory[38] <= 32'h0;
memory[39] <= 32'h0;
memory[40] <= 32'h0;
memory[41] <= 32'h0;
memory[42] <= 32'h0;
memory[43] <= 32'h0;
memory[44] <= 32'h0;
memory[45] <= 32'h0;
memory[46] <= 32'h0;
memory[47] <= 32'h0;
memory[48] <= 32'h0;
memory[49] <= 32'h0;
memory[50] <= 32'h0;
memory[51] <= 32'h0;
memory[52] <= 32'h0;
memory[53] <= 32'h0;
memory[54] <= 32'h0;
memory[55] <= 32'h0;
memory[56] <= 32'h0;
memory[57] <= 32'h0;
memory[58] <= 32'h0;
memory[59] <= 32'h0;
memory[60] <= 32'h0;
memory[61] <= 32'h0;
memory[62] <= 32'h1;
memory[63] <= 32'h1;
memory[64] <= 32'h1;
memory[65] <= 32'h1;
memory[66] <= 32'h0;
memory[67] <= 32'h0;
memory[68] <= 32'h0;
memory[69] <= 32'h0;
memory[70] <= 32'h0;
memory[71] <= 32'h0;
memory[72] <= 32'h0;
memory[73] <= 32'h0;
memory[74] <= 32'h0;
memory[75] <= 32'h0;
memory[76] <= 32'h0;
memory[77] <= 32'h0;
memory[78] <= 32'h0;
memory[79] <= 32'h0;
memory[80] <= 32'h0;
memory[81] <= 32'h0;
memory[82] <= 32'h0;
memory[83] <= 32'h0;
memory[84] <= 32'h0;
memory[85] <= 32'h0;
memory[86] <= 32'h0;
memory[87] <= 32'h0;
memory[88] <= 32'h0;
memory[89] <= 32'h0;
memory[90] <= 32'h0;
memory[91] <= 32'h0;
memory[92] <= 32'h0;
memory[93] <= 32'h1;
memory[94] <= 32'h1;
memory[95] <= 32'h1;
memory[96] <= 32'h1;
memory[97] <= 32'h0;
memory[98] <= 32'h0;
memory[99] <= 32'h0;
memory[100] <= 32'h0;
memory[101] <= 32'h0;
memory[102] <= 32'h0;
memory[103] <= 32'h0;
memory[104] <= 32'h0;
memory[105] <= 32'h0;
memory[106] <= 32'h0;
memory[107] <= 32'h0;
memory[108] <= 32'h0;
memory[109] <= 32'h0;
memory[110] <= 32'h0;
memory[111] <= 32'h0;
memory[112] <= 32'h0;
memory[113] <= 32'h0;
memory[114] <= 32'h0;
memory[115] <= 32'h0;
memory[116] <= 32'h0;
memory[117] <= 32'h0;
memory[118] <= 32'h0;
memory[119] <= 32'h0;
memory[120] <= 32'h0;
memory[121] <= 32'h0;
memory[122] <= 32'h0;
memory[123] <= 32'h0;
memory[124] <= 32'h1;
memory[125] <= 32'h1;
memory[126] <= 32'h1;
memory[127] <= 32'h1;
memory[128] <= 32'h0;
memory[129] <= 32'h0;
memory[130] <= 32'h0;
memory[131] <= 32'h0;
memory[132] <= 32'h0;
memory[133] <= 32'h0;
memory[134] <= 32'h0;
memory[135] <= 32'h0;
memory[136] <= 32'h0;
memory[137] <= 32'h0;
memory[138] <= 32'h0;
memory[139] <= 32'h0;
memory[140] <= 32'h0;
memory[141] <= 32'h0;
memory[142] <= 32'h0;
memory[143] <= 32'h0;
memory[144] <= 32'h0;
memory[145] <= 32'h0;
memory[146] <= 32'h0;
memory[147] <= 32'h0;
memory[148] <= 32'h0;
memory[149] <= 32'h0;
memory[150] <= 32'h0;
memory[151] <= 32'h0;
memory[152] <= 32'h0;
memory[153] <= 32'h0;
memory[154] <= 32'h0;
memory[155] <= 32'h1;
memory[156] <= 32'h1;
memory[157] <= 32'h1;
memory[158] <= 32'h1;
memory[159] <= 32'h0;
memory[160] <= 32'h0;
memory[161] <= 32'h0;
memory[162] <= 32'h0;
memory[163] <= 32'h0;
memory[164] <= 32'h0;
memory[165] <= 32'h0;
memory[166] <= 32'h0;
memory[167] <= 32'h0;
memory[168] <= 32'h0;
memory[169] <= 32'h0;
memory[170] <= 32'h0;
memory[171] <= 32'h0;
memory[172] <= 32'h0;
memory[173] <= 32'h0;
memory[174] <= 32'h0;
memory[175] <= 32'h0;
memory[176] <= 32'h0;
memory[177] <= 32'h0;
memory[178] <= 32'h0;
memory[179] <= 32'h0;
memory[180] <= 32'h0;
memory[181] <= 32'h0;
memory[182] <= 32'h0;
memory[183] <= 32'h0;
memory[184] <= 32'h0;
memory[185] <= 32'h0;
memory[186] <= 32'h1;
memory[187] <= 32'h1;
memory[188] <= 32'h1;
memory[189] <= 32'h1;
memory[190] <= 32'h0;
memory[191] <= 32'h0;
memory[192] <= 32'h0;
memory[193] <= 32'h0;
memory[194] <= 32'h0;
memory[195] <= 32'h0;
memory[196] <= 32'h0;
memory[197] <= 32'h0;
memory[198] <= 32'h0;
memory[199] <= 32'h0;
memory[200] <= 32'h0;
memory[201] <= 32'h0;
memory[202] <= 32'h0;
memory[203] <= 32'h0;
memory[204] <= 32'h0;
memory[205] <= 32'h0;
memory[206] <= 32'h0;
memory[207] <= 32'h0;
memory[208] <= 32'h0;
memory[209] <= 32'h0;
memory[210] <= 32'h0;
memory[211] <= 32'h0;
memory[212] <= 32'h0;
memory[213] <= 32'h0;
memory[214] <= 32'h0;
memory[215] <= 32'h0;
memory[216] <= 32'h0;
memory[217] <= 32'h1;
memory[218] <= 32'h1;
memory[219] <= 32'h1;
memory[220] <= 32'h1;
memory[221] <= 32'h0;
memory[222] <= 32'h0;
memory[223] <= 32'h0;
memory[224] <= 32'h0;
memory[225] <= 32'h0;
memory[226] <= 32'h0;
memory[227] <= 32'h0;
memory[228] <= 32'h0;
memory[229] <= 32'h0;
memory[230] <= 32'h0;
memory[231] <= 32'h0;
memory[232] <= 32'h0;
memory[233] <= 32'h0;
memory[234] <= 32'h0;
memory[235] <= 32'h0;
memory[236] <= 32'h0;
memory[237] <= 32'h0;
memory[238] <= 32'h0;
memory[239] <= 32'h0;
memory[240] <= 32'h0;
memory[241] <= 32'h0;
memory[242] <= 32'h0;
memory[243] <= 32'h0;
memory[244] <= 32'h0;
memory[245] <= 32'h0;
memory[246] <= 32'h0;
memory[247] <= 32'h0;
memory[248] <= 32'h1;
memory[249] <= 32'h1;
memory[250] <= 32'h1;
memory[251] <= 32'h1;
memory[252] <= 32'h0;
memory[253] <= 32'h0;
memory[254] <= 32'h0;
memory[255] <= 32'h0;
memory[256] <= 32'h0;
memory[257] <= 32'h0;
memory[258] <= 32'h0;
memory[259] <= 32'h0;
memory[260] <= 32'h0;
memory[261] <= 32'h0;
memory[262] <= 32'h0;
memory[263] <= 32'h0;
memory[264] <= 32'h0;
memory[265] <= 32'h0;
memory[266] <= 32'h0;
memory[267] <= 32'h0;
memory[268] <= 32'h0;
memory[269] <= 32'h0;
memory[270] <= 32'h0;
memory[271] <= 32'h0;
memory[272] <= 32'h0;
memory[273] <= 32'h0;
memory[274] <= 32'h0;
memory[275] <= 32'h0;
memory[276] <= 32'h0;
memory[277] <= 32'h0;
memory[278] <= 32'h0;
memory[279] <= 32'h0;
memory[280] <= 32'h0;
memory[281] <= 32'h0;
memory[282] <= 32'h0;
memory[283] <= 32'h0;
memory[284] <= 32'h0;
memory[285] <= 32'h0;
memory[286] <= 32'h0;
memory[287] <= 32'h0;
memory[288] <= 32'h0;
memory[289] <= 32'h0;
memory[290] <= 32'h0;
memory[291] <= 32'h0;
memory[292] <= 32'h0;
memory[293] <= 32'h0;
memory[294] <= 32'h0;
memory[295] <= 32'h0;
memory[296] <= 32'h0;
memory[297] <= 32'h0;
memory[298] <= 32'h0;
memory[299] <= 32'h0;
memory[300] <= 32'h0;
memory[301] <= 32'h0;
memory[302] <= 32'h0;
memory[303] <= 32'h0;
memory[304] <= 32'h0;
memory[305] <= 32'h0;
memory[306] <= 32'h0;
memory[307] <= 32'h0;
memory[308] <= 32'h0;
memory[309] <= 32'h0;
memory[310] <= 32'h0;
memory[311] <= 32'h0;
memory[312] <= 32'h0;
memory[313] <= 32'h0;
memory[314] <= 32'h0;
memory[315] <= 32'h0;
memory[316] <= 32'h0;
memory[317] <= 32'h0;
memory[318] <= 32'h0;
memory[319] <= 32'h0;
memory[320] <= 32'h0;
memory[321] <= 32'h0;
memory[322] <= 32'h0;
memory[323] <= 32'h0;
memory[324] <= 32'h0;
memory[325] <= 32'h0;
memory[326] <= 32'h0;
memory[327] <= 32'h0;
memory[328] <= 32'h0;
memory[329] <= 32'h0;
memory[330] <= 32'h0;
memory[331] <= 32'h0;
memory[332] <= 32'h0;
memory[333] <= 32'h0;
memory[334] <= 32'h0;
memory[335] <= 32'h0;
memory[336] <= 32'h0;
memory[337] <= 32'h0;
memory[338] <= 32'h0;
memory[339] <= 32'h0;
memory[340] <= 32'h0;
memory[341] <= 32'h0;
memory[342] <= 32'h0;
memory[343] <= 32'h0;
memory[344] <= 32'h0;
memory[345] <= 32'h0;
memory[346] <= 32'h0;
memory[347] <= 32'h0;
memory[348] <= 32'h0;
memory[349] <= 32'h0;
memory[350] <= 32'h0;
memory[351] <= 32'h0;
memory[352] <= 32'h0;
memory[353] <= 32'h0;
memory[354] <= 32'h0;
memory[355] <= 32'h0;
memory[356] <= 32'h0;
memory[357] <= 32'h0;
memory[358] <= 32'h0;
memory[359] <= 32'h0;
memory[360] <= 32'h0;
memory[361] <= 32'h0;
memory[362] <= 32'h0;
memory[363] <= 32'h0;
memory[364] <= 32'h0;
memory[365] <= 32'h0;
memory[366] <= 32'h0;
memory[367] <= 32'h0;
memory[368] <= 32'h0;
memory[369] <= 32'h0;
memory[370] <= 32'h0;
memory[371] <= 32'h0;
memory[372] <= 32'h0;
memory[373] <= 32'h0;
memory[374] <= 32'h0;
memory[375] <= 32'h0;
memory[376] <= 32'h0;
memory[377] <= 32'h0;
memory[378] <= 32'h0;
memory[379] <= 32'h0;
memory[380] <= 32'h0;
memory[381] <= 32'h0;
memory[382] <= 32'h0;
memory[383] <= 32'h0;
memory[384] <= 32'h0;
memory[385] <= 32'h0;
memory[386] <= 32'h0;
memory[387] <= 32'h0;
memory[388] <= 32'h0;
memory[389] <= 32'h0;
memory[390] <= 32'h0;
memory[391] <= 32'h0;
memory[392] <= 32'h0;
memory[393] <= 32'h0;
memory[394] <= 32'h0;
memory[395] <= 32'h0;
memory[396] <= 32'h0;
memory[397] <= 32'h0;
memory[398] <= 32'h0;
memory[399] <= 32'h0;
memory[400] <= 32'h0;
memory[401] <= 32'h0;
memory[402] <= 32'h0;
memory[403] <= 32'h0;
memory[404] <= 32'h0;
memory[405] <= 32'h0;
memory[406] <= 32'h0;
memory[407] <= 32'h0;
memory[408] <= 32'h0;
memory[409] <= 32'h0;
memory[410] <= 32'h0;
memory[411] <= 32'h0;
memory[412] <= 32'h0;
memory[413] <= 32'h0;
memory[414] <= 32'h0;
memory[415] <= 32'h0;
memory[416] <= 32'h0;
memory[417] <= 32'h0;
memory[418] <= 32'h0;
memory[419] <= 32'h0;
memory[420] <= 32'h0;
memory[421] <= 32'h0;
memory[422] <= 32'h0;
memory[423] <= 32'h0;
memory[424] <= 32'h0;
memory[425] <= 32'h0;
memory[426] <= 32'h0;
memory[427] <= 32'h0;
memory[428] <= 32'h0;
memory[429] <= 32'h0;
memory[430] <= 32'h0;
memory[431] <= 32'h0;
memory[432] <= 32'h0;
memory[433] <= 32'h0;
memory[434] <= 32'h0;
memory[435] <= 32'h0;
memory[436] <= 32'h0;
memory[437] <= 32'h0;
memory[438] <= 32'h0;
memory[439] <= 32'h0;
memory[440] <= 32'h0;
memory[441] <= 32'h0;
memory[442] <= 32'h0;
memory[443] <= 32'h0;
memory[444] <= 32'h0;
memory[445] <= 32'h0;
memory[446] <= 32'h0;
memory[447] <= 32'h0;
memory[448] <= 32'h0;
memory[449] <= 32'h0;
memory[450] <= 32'h0;
memory[451] <= 32'h0;
memory[452] <= 32'h0;
memory[453] <= 32'h0;
memory[454] <= 32'h0;
memory[455] <= 32'h0;
memory[456] <= 32'h0;
memory[457] <= 32'h0;
memory[458] <= 32'h0;
memory[459] <= 32'h0;
memory[460] <= 32'h0;
memory[461] <= 32'h0;
memory[462] <= 32'h0;
memory[463] <= 32'h0;
memory[464] <= 32'h0;
memory[465] <= 32'h0;
memory[466] <= 32'h0;
memory[467] <= 32'h0;
memory[468] <= 32'h0;
memory[469] <= 32'h0;
memory[470] <= 32'h0;
memory[471] <= 32'h0;
memory[472] <= 32'h0;
memory[473] <= 32'h0;
memory[474] <= 32'h0;
memory[475] <= 32'h0;
memory[476] <= 32'h0;
memory[477] <= 32'h0;
memory[478] <= 32'h0;
memory[479] <= 32'h0;
memory[480] <= 32'h0;
memory[481] <= 32'h0;
memory[482] <= 32'h0;
memory[483] <= 32'h0;
memory[484] <= 32'h0;
memory[485] <= 32'h0;
memory[486] <= 32'h0;
memory[487] <= 32'h0;
memory[488] <= 32'h0;
memory[489] <= 32'h0;
memory[490] <= 32'h0;
memory[491] <= 32'h0;
memory[492] <= 32'h0;
memory[493] <= 32'h0;
memory[494] <= 32'h0;
memory[495] <= 32'h0;
memory[496] <= 32'h0;
memory[497] <= 32'h0;
memory[498] <= 32'h0;
memory[499] <= 32'h0;
memory[500] <= 32'h0;
memory[501] <= 32'h0;
memory[502] <= 32'h0;
memory[503] <= 32'h0;
memory[504] <= 32'h0;
memory[505] <= 32'h0;
memory[506] <= 32'h0;
memory[507] <= 32'h0;
memory[508] <= 32'h0;
memory[509] <= 32'h0;
memory[510] <= 32'h0;
memory[511] <= 32'h0;
memory[512] <= 32'h0;
memory[513] <= 32'h0;
memory[514] <= 32'h0;
memory[515] <= 32'h0;
memory[516] <= 32'h0;
memory[517] <= 32'h0;
memory[518] <= 32'h0;
memory[519] <= 32'h0;
memory[520] <= 32'h0;
memory[521] <= 32'h0;
memory[522] <= 32'h0;
memory[523] <= 32'h0;
memory[524] <= 32'h0;
memory[525] <= 32'h0;
memory[526] <= 32'h0;
memory[527] <= 32'h0;
memory[528] <= 32'h0;
memory[529] <= 32'h0;
memory[530] <= 32'h0;
memory[531] <= 32'h0;
memory[532] <= 32'h0;
memory[533] <= 32'h0;
memory[534] <= 32'h0;
memory[535] <= 32'h0;
memory[536] <= 32'h0;
memory[537] <= 32'h0;
memory[538] <= 32'h0;
memory[539] <= 32'h0;
memory[540] <= 32'h0;
memory[541] <= 32'h0;
memory[542] <= 32'h0;
memory[543] <= 32'h0;
memory[544] <= 32'h0;
memory[545] <= 32'h0;
memory[546] <= 32'h0;
memory[547] <= 32'h0;
memory[548] <= 32'h0;
memory[549] <= 32'h0;
memory[550] <= 32'h0;
memory[551] <= 32'h0;
memory[552] <= 32'h0;
memory[553] <= 32'h0;
memory[554] <= 32'h0;
memory[555] <= 32'h0;
memory[556] <= 32'h0;
memory[557] <= 32'h0;
memory[558] <= 32'h0;
memory[559] <= 32'h0;
memory[560] <= 32'h0;
memory[561] <= 32'h0;
memory[562] <= 32'h0;
memory[563] <= 32'h0;
memory[564] <= 32'h0;
memory[565] <= 32'h0;
memory[566] <= 32'h0;
memory[567] <= 32'h0;
memory[568] <= 32'h0;
memory[569] <= 32'h0;
memory[570] <= 32'h0;
memory[571] <= 32'h0;
memory[572] <= 32'h0;
memory[573] <= 32'h0;
memory[574] <= 32'h0;
memory[575] <= 32'h0;
memory[576] <= 32'h0;
memory[577] <= 32'h0;
memory[578] <= 32'h0;
memory[579] <= 32'h0;
memory[580] <= 32'h0;
memory[581] <= 32'h0;
memory[582] <= 32'h0;
memory[583] <= 32'h0;
memory[584] <= 32'h0;
memory[585] <= 32'h0;
memory[586] <= 32'h0;
memory[587] <= 32'h0;
memory[588] <= 32'h0;
memory[589] <= 32'h0;
memory[590] <= 32'h0;
memory[591] <= 32'h0;
memory[592] <= 32'h0;
memory[593] <= 32'h0;
memory[594] <= 32'h0;
memory[595] <= 32'h0;
memory[596] <= 32'h0;
memory[597] <= 32'h0;
memory[598] <= 32'h0;
memory[599] <= 32'h0;
memory[600] <= 32'h0;
memory[601] <= 32'h0;
memory[602] <= 32'h0;
memory[603] <= 32'h0;
memory[604] <= 32'h0;
memory[605] <= 32'h0;
memory[606] <= 32'h0;
memory[607] <= 32'h0;
memory[608] <= 32'h0;
memory[609] <= 32'h0;
memory[610] <= 32'h0;
memory[611] <= 32'h0;
memory[612] <= 32'h0;
memory[613] <= 32'h0;
memory[614] <= 32'h0;
memory[615] <= 32'h0;
memory[616] <= 32'h0;
memory[617] <= 32'h0;
memory[618] <= 32'h0;
memory[619] <= 32'h0;
memory[620] <= 32'h0;
memory[621] <= 32'h0;
memory[622] <= 32'h0;
memory[623] <= 32'h0;
memory[624] <= 32'h0;
memory[625] <= 32'h0;
memory[626] <= 32'h0;
memory[627] <= 32'h0;
memory[628] <= 32'h0;
memory[629] <= 32'h0;
memory[630] <= 32'h0;
memory[631] <= 32'h0;
memory[632] <= 32'h0;
memory[633] <= 32'h0;
memory[634] <= 32'h0;
memory[635] <= 32'h0;
memory[636] <= 32'h0;
memory[637] <= 32'h0;
memory[638] <= 32'h0;
memory[639] <= 32'h0;
memory[640] <= 32'h0;
memory[641] <= 32'h0;
memory[642] <= 32'h0;
memory[643] <= 32'h0;
memory[644] <= 32'h0;
memory[645] <= 32'h0;
memory[646] <= 32'h0;
memory[647] <= 32'h0;
memory[648] <= 32'h0;
memory[649] <= 32'h0;
memory[650] <= 32'h0;
memory[651] <= 32'h0;
memory[652] <= 32'h0;
memory[653] <= 32'h0;
memory[654] <= 32'h0;
memory[655] <= 32'h0;
memory[656] <= 32'h0;
memory[657] <= 32'h0;
memory[658] <= 32'h0;
memory[659] <= 32'h0;
memory[660] <= 32'h0;
memory[661] <= 32'h0;
memory[662] <= 32'h0;
memory[663] <= 32'h0;
memory[664] <= 32'h0;
memory[665] <= 32'h0;
memory[666] <= 32'h0;
memory[667] <= 32'h0;
memory[668] <= 32'h0;
memory[669] <= 32'h0;
memory[670] <= 32'h0;
memory[671] <= 32'h0;
memory[672] <= 32'h0;
memory[673] <= 32'h0;
memory[674] <= 32'h0;
memory[675] <= 32'h0;
memory[676] <= 32'h0;
memory[677] <= 32'h0;
memory[678] <= 32'h0;
memory[679] <= 32'h0;
memory[680] <= 32'h0;
memory[681] <= 32'h0;
memory[682] <= 32'h0;
memory[683] <= 32'h0;
memory[684] <= 32'h0;
memory[685] <= 32'h0;
memory[686] <= 32'h0;
memory[687] <= 32'h0;
memory[688] <= 32'h0;
memory[689] <= 32'h0;
memory[690] <= 32'h0;
memory[691] <= 32'h0;
memory[692] <= 32'h0;
memory[693] <= 32'h0;
memory[694] <= 32'h0;
memory[695] <= 32'h0;
memory[696] <= 32'h0;
memory[697] <= 32'h0;
memory[698] <= 32'h0;
memory[699] <= 32'h0;
memory[700] <= 32'h0;
memory[701] <= 32'h0;
memory[702] <= 32'h0;
memory[703] <= 32'h0;
memory[704] <= 32'h0;
memory[705] <= 32'h0;
memory[706] <= 32'h0;
memory[707] <= 32'h0;
memory[708] <= 32'h0;
memory[709] <= 32'h0;
memory[710] <= 32'h0;
memory[711] <= 32'h0;
memory[712] <= 32'h0;
memory[713] <= 32'h0;
memory[714] <= 32'h0;
memory[715] <= 32'h0;
memory[716] <= 32'h0;
memory[717] <= 32'h0;
memory[718] <= 32'h0;
memory[719] <= 32'h0;
memory[720] <= 32'h0;
memory[721] <= 32'h0;
memory[722] <= 32'h0;
memory[723] <= 32'h0;
memory[724] <= 32'h0;
memory[725] <= 32'h0;
memory[726] <= 32'h0;
memory[727] <= 32'h0;
memory[728] <= 32'h0;
memory[729] <= 32'h0;
memory[730] <= 32'h0;
memory[731] <= 32'h0;
memory[732] <= 32'h0;
memory[733] <= 32'h0;
memory[734] <= 32'h0;
memory[735] <= 32'h0;
memory[736] <= 32'h0;
memory[737] <= 32'h0;
memory[738] <= 32'h0;
memory[739] <= 32'h0;
memory[740] <= 32'h0;
memory[741] <= 32'h0;
memory[742] <= 32'h0;
memory[743] <= 32'h0;
memory[744] <= 32'h0;
memory[745] <= 32'h0;
memory[746] <= 32'h0;
memory[747] <= 32'h0;
memory[748] <= 32'h0;
memory[749] <= 32'h0;
memory[750] <= 32'h0;
memory[751] <= 32'h0;
memory[752] <= 32'h0;
memory[753] <= 32'h0;
memory[754] <= 32'h0;
memory[755] <= 32'h0;
memory[756] <= 32'h0;
memory[757] <= 32'h0;
memory[758] <= 32'h0;
memory[759] <= 32'h0;
memory[760] <= 32'h0;
memory[761] <= 32'h0;
memory[762] <= 32'h0;
memory[763] <= 32'h0;
memory[764] <= 32'h0;
memory[765] <= 32'h0;
memory[766] <= 32'h0;
memory[767] <= 32'h0;
memory[768] <= 32'h0;
memory[769] <= 32'h0;
memory[770] <= 32'h0;
memory[771] <= 32'h0;
memory[772] <= 32'h0;
memory[773] <= 32'h0;
memory[774] <= 32'h0;
memory[775] <= 32'h0;
memory[776] <= 32'h0;
memory[777] <= 32'h0;
memory[778] <= 32'h0;
memory[779] <= 32'h0;
memory[780] <= 32'h0;
memory[781] <= 32'h0;
memory[782] <= 32'h0;
memory[783] <= 32'h0;
memory[784] <= 32'h0;
memory[785] <= 32'h0;
memory[786] <= 32'h0;
memory[787] <= 32'h0;
memory[788] <= 32'h0;
memory[789] <= 32'h0;
memory[790] <= 32'h0;
memory[791] <= 32'h0;
memory[792] <= 32'h0;
memory[793] <= 32'h0;
memory[794] <= 32'h0;
memory[795] <= 32'h0;
memory[796] <= 32'h0;
memory[797] <= 32'h0;
memory[798] <= 32'h0;
memory[799] <= 32'h0;
memory[800] <= 32'h0;
memory[801] <= 32'h0;
memory[802] <= 32'h0;
memory[803] <= 32'h0;
memory[804] <= 32'h0;
memory[805] <= 32'h0;
memory[806] <= 32'h0;
memory[807] <= 32'h0;
memory[808] <= 32'h0;
memory[809] <= 32'h0;
memory[810] <= 32'h0;
memory[811] <= 32'h0;
memory[812] <= 32'h0;
memory[813] <= 32'h0;
memory[814] <= 32'h0;
memory[815] <= 32'h0;
memory[816] <= 32'h0;
memory[817] <= 32'h0;
memory[818] <= 32'h0;
memory[819] <= 32'h0;
memory[820] <= 32'h0;
memory[821] <= 32'h0;
memory[822] <= 32'h0;
memory[823] <= 32'h0;
memory[824] <= 32'h0;
memory[825] <= 32'h0;
memory[826] <= 32'h0;
memory[827] <= 32'h0;
memory[828] <= 32'h0;
memory[829] <= 32'h0;
memory[830] <= 32'h0;
memory[831] <= 32'h0;
memory[832] <= 32'h0;
memory[833] <= 32'h0;
memory[834] <= 32'h0;
memory[835] <= 32'h0;
memory[836] <= 32'h0;
memory[837] <= 32'h0;
memory[838] <= 32'h0;
memory[839] <= 32'h0;
memory[840] <= 32'h0;
memory[841] <= 32'h0;
memory[842] <= 32'h0;
memory[843] <= 32'h0;
memory[844] <= 32'h0;
memory[845] <= 32'h0;
memory[846] <= 32'h0;
memory[847] <= 32'h0;
memory[848] <= 32'h0;
memory[849] <= 32'h0;
memory[850] <= 32'h0;
memory[851] <= 32'h0;
memory[852] <= 32'h0;
memory[853] <= 32'h0;
memory[854] <= 32'h0;
memory[855] <= 32'h0;
memory[856] <= 32'h0;
memory[857] <= 32'h0;
memory[858] <= 32'h0;
memory[859] <= 32'h0;
memory[860] <= 32'h0;
memory[861] <= 32'h0;
memory[862] <= 32'h0;
memory[863] <= 32'h0;
memory[864] <= 32'h0;
memory[865] <= 32'h0;
memory[866] <= 32'h0;
memory[867] <= 32'h0;
memory[868] <= 32'h0;
memory[869] <= 32'h0;
memory[870] <= 32'h0;
memory[871] <= 32'h0;
memory[872] <= 32'h0;
memory[873] <= 32'h0;
memory[874] <= 32'h0;
memory[875] <= 32'h0;
memory[876] <= 32'h0;
memory[877] <= 32'h0;
memory[878] <= 32'h0;
memory[879] <= 32'h0;
memory[880] <= 32'h0;
memory[881] <= 32'h0;
memory[882] <= 32'h0;
memory[883] <= 32'h0;
memory[884] <= 32'h0;
memory[885] <= 32'h0;
memory[886] <= 32'h0;
memory[887] <= 32'h0;
memory[888] <= 32'h0;
memory[889] <= 32'h0;
memory[890] <= 32'h0;
memory[891] <= 32'h0;
memory[892] <= 32'h0;
memory[893] <= 32'h0;
memory[894] <= 32'h0;
memory[895] <= 32'h0;
memory[896] <= 32'h0;
memory[897] <= 32'h0;
memory[898] <= 32'h0;
memory[899] <= 32'h0;
memory[900] <= 32'h0;
memory[901] <= 32'h0;
memory[902] <= 32'h0;
memory[903] <= 32'h0;
memory[904] <= 32'h0;
memory[905] <= 32'h0;
memory[906] <= 32'h0;
memory[907] <= 32'h0;
memory[908] <= 32'h0;
memory[909] <= 32'h0;
memory[910] <= 32'h0;
memory[911] <= 32'h0;
memory[912] <= 32'h0;
memory[913] <= 32'h0;
memory[914] <= 32'h0;
memory[915] <= 32'h0;
memory[916] <= 32'h0;
memory[917] <= 32'h0;
memory[918] <= 32'h0;
memory[919] <= 32'h0;
memory[920] <= 32'h0;
memory[921] <= 32'h0;
memory[922] <= 32'h0;
memory[923] <= 32'h0;
memory[924] <= 32'h0;
memory[925] <= 32'h0;
memory[926] <= 32'h0;
memory[927] <= 32'h0;
memory[928] <= 32'h0;
memory[929] <= 32'h0;
memory[930] <= 32'h0;
memory[931] <= 32'h0;
memory[932] <= 32'h0;
memory[933] <= 32'h0;
memory[934] <= 32'h0;
memory[935] <= 32'h0;
memory[936] <= 32'h0;
memory[937] <= 32'h0;
memory[938] <= 32'h0;
memory[939] <= 32'h0;
memory[940] <= 32'h0;
memory[941] <= 32'h0;
memory[942] <= 32'h0;
memory[943] <= 32'h0;
memory[944] <= 32'h0;
memory[945] <= 32'h0;
memory[946] <= 32'h0;
memory[947] <= 32'h0;
memory[948] <= 32'h0;
memory[949] <= 32'h0;
memory[950] <= 32'h0;
memory[951] <= 32'h0;
memory[952] <= 32'h0;
memory[953] <= 32'h0;
memory[954] <= 32'h0;
memory[955] <= 32'h0;
memory[956] <= 32'h0;
memory[957] <= 32'h0;
memory[958] <= 32'h0;
memory[959] <= 32'h0;
memory[960] <= 32'h0;
memory[961] <= 32'h0;
memory[962] <= 32'h0;
memory[963] <= 32'h0;
memory[964] <= 32'h0;
memory[965] <= 32'h0;
memory[966] <= 32'h0;
memory[967] <= 32'h0;
memory[968] <= 32'h0;
memory[969] <= 32'h0;
memory[970] <= 32'h0;
memory[971] <= 32'h0;
memory[972] <= 32'h0;
memory[973] <= 32'h0;
memory[974] <= 32'h0;
memory[975] <= 32'h0;
memory[976] <= 32'h0;
memory[977] <= 32'h0;
memory[978] <= 32'h0;
memory[979] <= 32'h0;
memory[980] <= 32'h0;
memory[981] <= 32'h0;
memory[982] <= 32'h0;
memory[983] <= 32'h0;
memory[984] <= 32'h0;
memory[985] <= 32'h0;
memory[986] <= 32'h0;
memory[987] <= 32'h0;
memory[988] <= 32'h0;
memory[989] <= 32'h0;
memory[990] <= 32'h0;
memory[991] <= 32'h0;
memory[992] <= 32'h0;
memory[993] <= 32'h0;
memory[994] <= 32'h0;
memory[995] <= 32'h0;
memory[996] <= 32'h0;
memory[997] <= 32'h0;
memory[998] <= 32'h0;
memory[999] <= 32'h0;
memory[1000] <= 32'h0;
memory[1001] <= 32'h0;
memory[1002] <= 32'h0;
memory[1003] <= 32'h0;
memory[1004] <= 32'h0;
memory[1005] <= 32'h0;
memory[1006] <= 32'h0;
memory[1007] <= 32'h0;
memory[1008] <= 32'h0;
memory[1009] <= 32'h0;
memory[1010] <= 32'h0;
memory[1011] <= 32'h0;
memory[1012] <= 32'h0;
memory[1013] <= 32'h0;
memory[1014] <= 32'h0;
memory[1015] <= 32'h0;
memory[1016] <= 32'h0;
memory[1017] <= 32'h0;
memory[1018] <= 32'h0;
memory[1019] <= 32'h0;
memory[1020] <= 32'h0;
memory[1021] <= 32'h0;
memory[1022] <= 32'h0;
memory[1023] <= 32'h0;
memory[1024] <= 32'h0;
memory[1025] <= 32'h0;
memory[1026] <= 32'h0;
memory[1027] <= 32'h0;
memory[1028] <= 32'h0;
memory[1029] <= 32'h0;
memory[1030] <= 32'h0;
memory[1031] <= 32'h0;
memory[1032] <= 32'h0;
memory[1033] <= 32'h0;
memory[1034] <= 32'h0;
memory[1035] <= 32'h0;
memory[1036] <= 32'h0;
memory[1037] <= 32'h0;
memory[1038] <= 32'h0;
memory[1039] <= 32'h0;
memory[1040] <= 32'h0;
memory[1041] <= 32'h0;
memory[1042] <= 32'h0;
memory[1043] <= 32'h0;
memory[1044] <= 32'h0;
memory[1045] <= 32'h0;
memory[1046] <= 32'h0;
memory[1047] <= 32'h0;
memory[1048] <= 32'h0;
memory[1049] <= 32'h0;
memory[1050] <= 32'h0;
memory[1051] <= 32'h0;
memory[1052] <= 32'h0;
memory[1053] <= 32'h0;
memory[1054] <= 32'h0;
memory[1055] <= 32'h0;
memory[1056] <= 32'h0;
memory[1057] <= 32'h0;
memory[1058] <= 32'h0;
memory[1059] <= 32'h0;
memory[1060] <= 32'h0;
memory[1061] <= 32'h0;
memory[1062] <= 32'h0;
memory[1063] <= 32'h0;
memory[1064] <= 32'h0;
memory[1065] <= 32'h0;
memory[1066] <= 32'h0;
memory[1067] <= 32'h0;
memory[1068] <= 32'h0;
memory[1069] <= 32'h0;
memory[1070] <= 32'h0;
memory[1071] <= 32'h0;
memory[1072] <= 32'h0;
memory[1073] <= 32'h0;
memory[1074] <= 32'h0;
memory[1075] <= 32'h0;
memory[1076] <= 32'h0;
memory[1077] <= 32'h0;
memory[1078] <= 32'h0;
memory[1079] <= 32'h0;
memory[1080] <= 32'h0;
memory[1081] <= 32'h0;
memory[1082] <= 32'h0;
memory[1083] <= 32'h0;
memory[1084] <= 32'h0;
memory[1085] <= 32'h0;
memory[1086] <= 32'h0;
memory[1087] <= 32'h0;
memory[1088] <= 32'h0;
memory[1089] <= 32'h0;
memory[1090] <= 32'h0;
memory[1091] <= 32'h0;
memory[1092] <= 32'h0;
memory[1093] <= 32'h0;
memory[1094] <= 32'h0;
memory[1095] <= 32'h0;
memory[1096] <= 32'h0;
memory[1097] <= 32'h0;
memory[1098] <= 32'h0;
memory[1099] <= 32'h0;
memory[1100] <= 32'h0;
memory[1101] <= 32'h0;
memory[1102] <= 32'h0;
memory[1103] <= 32'h0;
memory[1104] <= 32'h0;
memory[1105] <= 32'h0;
memory[1106] <= 32'h0;
memory[1107] <= 32'h0;
memory[1108] <= 32'h0;
memory[1109] <= 32'h0;
memory[1110] <= 32'h0;
memory[1111] <= 32'h0;
memory[1112] <= 32'h0;
memory[1113] <= 32'h0;
memory[1114] <= 32'h0;
memory[1115] <= 32'h0;
memory[1116] <= 32'h0;
memory[1117] <= 32'h0;
memory[1118] <= 32'h0;
memory[1119] <= 32'h0;
memory[1120] <= 32'h0;
memory[1121] <= 32'h0;
memory[1122] <= 32'h0;
memory[1123] <= 32'h0;
memory[1124] <= 32'h0;
memory[1125] <= 32'h0;
memory[1126] <= 32'h0;
memory[1127] <= 32'h0;
memory[1128] <= 32'h0;
memory[1129] <= 32'h0;
memory[1130] <= 32'h0;
memory[1131] <= 32'h0;
memory[1132] <= 32'h0;
memory[1133] <= 32'h0;
memory[1134] <= 32'h0;
memory[1135] <= 32'h0;
memory[1136] <= 32'h0;
memory[1137] <= 32'h0;
memory[1138] <= 32'h0;
memory[1139] <= 32'h0;
memory[1140] <= 32'h0;
memory[1141] <= 32'h0;
memory[1142] <= 32'h0;
memory[1143] <= 32'h0;
memory[1144] <= 32'h0;
memory[1145] <= 32'h0;
memory[1146] <= 32'h0;
memory[1147] <= 32'h0;
memory[1148] <= 32'h0;
memory[1149] <= 32'h0;
memory[1150] <= 32'h0;
memory[1151] <= 32'h0;
memory[1152] <= 32'h0;
memory[1153] <= 32'h0;
memory[1154] <= 32'h0;
memory[1155] <= 32'h0;
memory[1156] <= 32'h0;
memory[1157] <= 32'h0;
memory[1158] <= 32'h0;
memory[1159] <= 32'h0;
memory[1160] <= 32'h0;
memory[1161] <= 32'h0;
memory[1162] <= 32'h0;
memory[1163] <= 32'h0;
memory[1164] <= 32'h0;
memory[1165] <= 32'h0;
memory[1166] <= 32'h0;
memory[1167] <= 32'h0;
memory[1168] <= 32'h0;
memory[1169] <= 32'h0;
memory[1170] <= 32'h0;
memory[1171] <= 32'h0;
memory[1172] <= 32'h0;
memory[1173] <= 32'h0;
memory[1174] <= 32'h0;
memory[1175] <= 32'h0;
memory[1176] <= 32'h0;
memory[1177] <= 32'h0;
memory[1178] <= 32'h0;
memory[1179] <= 32'h0;
memory[1180] <= 32'h0;
memory[1181] <= 32'h0;
memory[1182] <= 32'h0;
memory[1183] <= 32'h0;
memory[1184] <= 32'h0;
memory[1185] <= 32'h0;
memory[1186] <= 32'h0;
memory[1187] <= 32'h0;
memory[1188] <= 32'h0;
memory[1189] <= 32'h0;
memory[1190] <= 32'h0;
memory[1191] <= 32'h0;
memory[1192] <= 32'h0;
memory[1193] <= 32'h0;
memory[1194] <= 32'h0;
memory[1195] <= 32'h0;
memory[1196] <= 32'h0;
memory[1197] <= 32'h0;
memory[1198] <= 32'h0;
memory[1199] <= 32'h0;
memory[1200] <= 32'h0;
memory[1201] <= 32'h0;
memory[1202] <= 32'h0;
memory[1203] <= 32'h0;
memory[1204] <= 32'h0;
memory[1205] <= 32'h0;
memory[1206] <= 32'h0;
memory[1207] <= 32'h0;
memory[1208] <= 32'h0;
memory[1209] <= 32'h0;
memory[1210] <= 32'h0;
memory[1211] <= 32'h0;
memory[1212] <= 32'h0;
memory[1213] <= 32'h1;
memory[1214] <= 32'h1;
memory[1215] <= 32'h1;
memory[1216] <= 32'h1;
memory[1217] <= 32'h1;
memory[1218] <= 32'h1;
memory[1219] <= 32'h1;
memory[1220] <= 32'h1;
memory[1221] <= 32'h1;
memory[1222] <= 32'h1;
memory[1223] <= 32'h1;
memory[1224] <= 32'h1;
memory[1225] <= 32'h1;
memory[1226] <= 32'h1;
memory[1227] <= 32'h1;
memory[1228] <= 32'h1;
memory[1229] <= 32'h1;
memory[1230] <= 32'h1;
memory[1231] <= 32'h1;
memory[1232] <= 32'h1;
memory[1233] <= 32'h1;
memory[1234] <= 32'h1;
memory[1235] <= 32'h1;
memory[1236] <= 32'h1;
memory[1237] <= 32'h1;
memory[1238] <= 32'h1;
memory[1239] <= 32'h1;
memory[1240] <= 32'h1;
memory[1241] <= 32'h1;
memory[1242] <= 32'h1;
memory[1243] <= 32'h1;
memory[1244] <= 32'h1;
memory[1245] <= 32'h32;
memory[1246] <= 32'h1f;
memory[1247] <= 32'h8;
memory[1248] <= 32'h4;
memory[1249] <= 32'h0;
memory[1250] <= 32'h0;
memory[1251] <= 32'h0;
memory[1252] <= 32'h0;
memory[1253] <= 32'h0;
memory[1254] <= 32'h0;
memory[1255] <= 32'h0;
memory[1256] <= 32'h0;
memory[1257] <= 32'h0;
memory[1258] <= 32'h0;
memory[1259] <= 32'h0;
memory[1260] <= 32'h0;
memory[1261] <= 32'h0;
memory[1262] <= 32'h0;
memory[1263] <= 32'h0;
memory[1264] <= 32'h0;
memory[1265] <= 32'h0;
memory[1266] <= 32'h0;
memory[1267] <= 32'h0;
memory[1268] <= 32'h0;
memory[1269] <= 32'h0;
memory[1270] <= 32'h0;
memory[1271] <= 32'h0;
memory[1272] <= 32'h0;
memory[1273] <= 32'h0;
memory[1274] <= 32'h0;
memory[1275] <= 32'h0;
memory[1276] <= 32'h0;
memory[1277] <= 32'h0;
memory[1278] <= 32'h0;
memory[1279] <= 32'h0;
memory[1280] <= 32'h0;
memory[1281] <= 32'h0;
memory[1282] <= 32'h0;
memory[1283] <= 32'h0;
memory[1284] <= 32'h0;
memory[1285] <= 32'h0;
memory[1286] <= 32'h0;
memory[1287] <= 32'h0;
memory[1288] <= 32'h0;
memory[1289] <= 32'h0;
memory[1290] <= 32'h0;
memory[1291] <= 32'h0;
memory[1292] <= 32'h0;
memory[1293] <= 32'h0;
memory[1294] <= 32'h0;
memory[1295] <= 32'h0;
memory[1296] <= 32'h0;
memory[1297] <= 32'h0;
memory[1298] <= 32'h0;
memory[1299] <= 32'h0;
memory[1300] <= 32'h0;
memory[1301] <= 32'h0;
memory[1302] <= 32'h0;
memory[1303] <= 32'h0;
memory[1304] <= 32'h0;
memory[1305] <= 32'h0;
memory[1306] <= 32'h0;
memory[1307] <= 32'h0;
memory[1308] <= 32'h0;
memory[1309] <= 32'h0;
memory[1310] <= 32'h0;
memory[1311] <= 32'h0;
memory[1312] <= 32'h0;
memory[1313] <= 32'h0;
memory[1314] <= 32'h0;
memory[1315] <= 32'h0;
memory[1316] <= 32'h0;
memory[1317] <= 32'h0;
memory[1318] <= 32'h0;
memory[1319] <= 32'h0;
memory[1320] <= 32'h0;
memory[1321] <= 32'h0;
memory[1322] <= 32'h0;
memory[1323] <= 32'h0;
memory[1324] <= 32'h0;
memory[1325] <= 32'h0;
memory[1326] <= 32'h0;
memory[1327] <= 32'h0;
memory[1328] <= 32'h0;
memory[1329] <= 32'h0;
memory[1330] <= 32'h0;
memory[1331] <= 32'h0;
memory[1332] <= 32'h0;
memory[1333] <= 32'h0;
memory[1334] <= 32'h0;
memory[1335] <= 32'h0;
memory[1336] <= 32'h0;
memory[1337] <= 32'h0;
memory[1338] <= 32'h0;
memory[1339] <= 32'h0;
memory[1340] <= 32'h0;
memory[1341] <= 32'h0;
memory[1342] <= 32'h0;
memory[1343] <= 32'h0;
memory[1344] <= 32'h0;
memory[1345] <= 32'h0;
memory[1346] <= 32'h0;
memory[1347] <= 32'h0;
memory[1348] <= 32'h0;
memory[1349] <= 32'h0;
memory[1350] <= 32'h0;
memory[1351] <= 32'h0;
memory[1352] <= 32'h0;
memory[1353] <= 32'h0;
memory[1354] <= 32'h0;
memory[1355] <= 32'h0;
memory[1356] <= 32'h0;
memory[1357] <= 32'h0;
memory[1358] <= 32'h0;
memory[1359] <= 32'h0;
memory[1360] <= 32'h0;
memory[1361] <= 32'h0;
memory[1362] <= 32'h0;
memory[1363] <= 32'h0;
memory[1364] <= 32'h0;
memory[1365] <= 32'h0;
memory[1366] <= 32'h0;
memory[1367] <= 32'h0;
memory[1368] <= 32'h0;
memory[1369] <= 32'h0;
memory[1370] <= 32'h0;
memory[1371] <= 32'h0;
memory[1372] <= 32'h0;
memory[1373] <= 32'h0;
memory[1374] <= 32'h0;
memory[1375] <= 32'h0;
memory[1376] <= 32'h0;
memory[1377] <= 32'h0;
memory[1378] <= 32'h0;
memory[1379] <= 32'h0;
memory[1380] <= 32'h0;
memory[1381] <= 32'h0;
memory[1382] <= 32'h0;
memory[1383] <= 32'h0;
memory[1384] <= 32'h0;
memory[1385] <= 32'h0;
memory[1386] <= 32'h0;
memory[1387] <= 32'h0;
memory[1388] <= 32'h0;
memory[1389] <= 32'h0;
memory[1390] <= 32'h0;
memory[1391] <= 32'h0;
memory[1392] <= 32'h0;
memory[1393] <= 32'h0;
memory[1394] <= 32'h0;
memory[1395] <= 32'h0;
memory[1396] <= 32'h0;
memory[1397] <= 32'h0;
memory[1398] <= 32'h0;
memory[1399] <= 32'h0;
memory[1400] <= 32'h0;
memory[1401] <= 32'h0;
memory[1402] <= 32'h0;
memory[1403] <= 32'h0;
memory[1404] <= 32'h0;
memory[1405] <= 32'h0;
memory[1406] <= 32'h0;
memory[1407] <= 32'h0;
memory[1408] <= 32'h0;
memory[1409] <= 32'h0;
memory[1410] <= 32'h0;
memory[1411] <= 32'h0;
memory[1412] <= 32'h0;
memory[1413] <= 32'h0;
memory[1414] <= 32'h0;
memory[1415] <= 32'h0;
memory[1416] <= 32'h0;
memory[1417] <= 32'h0;
memory[1418] <= 32'h0;
memory[1419] <= 32'h0;
memory[1420] <= 32'h0;
memory[1421] <= 32'h0;
memory[1422] <= 32'h0;
memory[1423] <= 32'h0;
memory[1424] <= 32'h0;
memory[1425] <= 32'h0;
memory[1426] <= 32'h0;
memory[1427] <= 32'h0;
memory[1428] <= 32'h0;
memory[1429] <= 32'h0;
memory[1430] <= 32'h0;
memory[1431] <= 32'h0;
memory[1432] <= 32'h0;
memory[1433] <= 32'h0;
memory[1434] <= 32'h0;
memory[1435] <= 32'h0;
memory[1436] <= 32'h0;
memory[1437] <= 32'h0;
memory[1438] <= 32'h0;
memory[1439] <= 32'h0;
memory[1440] <= 32'h0;
memory[1441] <= 32'h0;
memory[1442] <= 32'h0;
memory[1443] <= 32'h0;
memory[1444] <= 32'h0;
memory[1445] <= 32'h0;
memory[1446] <= 32'h0;
memory[1447] <= 32'h0;
memory[1448] <= 32'h0;
memory[1449] <= 32'h0;
memory[1450] <= 32'h0;
memory[1451] <= 32'h0;
memory[1452] <= 32'h0;
memory[1453] <= 32'h0;
memory[1454] <= 32'h0;
memory[1455] <= 32'h0;
memory[1456] <= 32'h0;
memory[1457] <= 32'h0;
memory[1458] <= 32'h0;
memory[1459] <= 32'h0;
memory[1460] <= 32'h0;
memory[1461] <= 32'h0;
memory[1462] <= 32'h0;
memory[1463] <= 32'h0;
memory[1464] <= 32'h0;
memory[1465] <= 32'h0;
memory[1466] <= 32'h0;
memory[1467] <= 32'h0;
memory[1468] <= 32'h0;
memory[1469] <= 32'h0;
memory[1470] <= 32'h0;
memory[1471] <= 32'h0;
memory[1472] <= 32'h0;
memory[1473] <= 32'h0;
memory[1474] <= 32'h0;
memory[1475] <= 32'h0;
memory[1476] <= 32'h0;
memory[1477] <= 32'h0;
memory[1478] <= 32'h0;
memory[1479] <= 32'h0;
memory[1480] <= 32'h0;
memory[1481] <= 32'h0;
memory[1482] <= 32'h0;
memory[1483] <= 32'h0;
memory[1484] <= 32'h0;
memory[1485] <= 32'h0;
memory[1486] <= 32'h0;
memory[1487] <= 32'h0;
memory[1488] <= 32'h0;
memory[1489] <= 32'h0;
memory[1490] <= 32'h0;
memory[1491] <= 32'h0;
memory[1492] <= 32'h0;
memory[1493] <= 32'h0;
memory[1494] <= 32'h0;
memory[1495] <= 32'h0;
memory[1496] <= 32'h0;
memory[1497] <= 32'h0;
memory[1498] <= 32'h0;
memory[1499] <= 32'h0;
memory[1500] <= 32'h0;
memory[1501] <= 32'h0;
memory[1502] <= 32'h0;
memory[1503] <= 32'h0;
memory[1504] <= 32'h0;
memory[1505] <= 32'h0;
memory[1506] <= 32'h0;
memory[1507] <= 32'h0;
memory[1508] <= 32'h0;
memory[1509] <= 32'h0;
memory[1510] <= 32'h0;
memory[1511] <= 32'h0;
memory[1512] <= 32'h0;
memory[1513] <= 32'h0;
memory[1514] <= 32'h0;
memory[1515] <= 32'h0;
memory[1516] <= 32'h0;
memory[1517] <= 32'h0;
memory[1518] <= 32'h0;
memory[1519] <= 32'h0;
memory[1520] <= 32'h0;
memory[1521] <= 32'h0;
memory[1522] <= 32'h0;
memory[1523] <= 32'h0;
memory[1524] <= 32'h0;
memory[1525] <= 32'h0;
memory[1526] <= 32'h0;
memory[1527] <= 32'h0;
memory[1528] <= 32'h0;
memory[1529] <= 32'h0;
memory[1530] <= 32'h0;
memory[1531] <= 32'h0;
memory[1532] <= 32'h0;
memory[1533] <= 32'h0;
memory[1534] <= 32'h0;
memory[1535] <= 32'h0;
memory[1536] <= 32'h0;
memory[1537] <= 32'h0;
memory[1538] <= 32'h0;
memory[1539] <= 32'h0;
memory[1540] <= 32'h0;
memory[1541] <= 32'h0;
memory[1542] <= 32'h0;
memory[1543] <= 32'h0;
memory[1544] <= 32'h0;
memory[1545] <= 32'h0;
memory[1546] <= 32'h0;
memory[1547] <= 32'h0;
memory[1548] <= 32'h0;
memory[1549] <= 32'h0;
memory[1550] <= 32'h0;
memory[1551] <= 32'h0;
memory[1552] <= 32'h0;
memory[1553] <= 32'h0;
memory[1554] <= 32'h0;
memory[1555] <= 32'h0;
memory[1556] <= 32'h0;
memory[1557] <= 32'h0;
memory[1558] <= 32'h0;
memory[1559] <= 32'h0;
memory[1560] <= 32'h0;
memory[1561] <= 32'h0;
memory[1562] <= 32'h0;
memory[1563] <= 32'h0;
memory[1564] <= 32'h0;
memory[1565] <= 32'h0;
memory[1566] <= 32'h0;
memory[1567] <= 32'h0;
memory[1568] <= 32'h0;
memory[1569] <= 32'h0;
memory[1570] <= 32'h0;
memory[1571] <= 32'h0;
memory[1572] <= 32'h0;
memory[1573] <= 32'h0;
memory[1574] <= 32'h0;
memory[1575] <= 32'h0;
memory[1576] <= 32'h0;
memory[1577] <= 32'h0;
memory[1578] <= 32'h0;
memory[1579] <= 32'h0;
memory[1580] <= 32'h0;
memory[1581] <= 32'h0;
memory[1582] <= 32'h0;
memory[1583] <= 32'h0;
memory[1584] <= 32'h0;
memory[1585] <= 32'h0;
memory[1586] <= 32'h0;
memory[1587] <= 32'h0;
memory[1588] <= 32'h0;
memory[1589] <= 32'h0;
memory[1590] <= 32'h0;
memory[1591] <= 32'h0;
memory[1592] <= 32'h0;
memory[1593] <= 32'h0;
memory[1594] <= 32'h0;
memory[1595] <= 32'h0;
memory[1596] <= 32'h0;
memory[1597] <= 32'h0;
memory[1598] <= 32'h0;
memory[1599] <= 32'h0;
memory[1600] <= 32'h0;
memory[1601] <= 32'h0;
memory[1602] <= 32'h0;
memory[1603] <= 32'h0;
memory[1604] <= 32'h0;
memory[1605] <= 32'h0;
memory[1606] <= 32'h0;
memory[1607] <= 32'h0;
memory[1608] <= 32'h0;
memory[1609] <= 32'h0;
memory[1610] <= 32'h0;
memory[1611] <= 32'h0;
memory[1612] <= 32'h0;
memory[1613] <= 32'h0;
memory[1614] <= 32'h0;
memory[1615] <= 32'h0;
memory[1616] <= 32'h0;
memory[1617] <= 32'h0;
memory[1618] <= 32'h0;
memory[1619] <= 32'h0;
memory[1620] <= 32'h0;
memory[1621] <= 32'h0;
memory[1622] <= 32'h0;
memory[1623] <= 32'h0;
memory[1624] <= 32'h0;
memory[1625] <= 32'h0;
memory[1626] <= 32'h0;
memory[1627] <= 32'h0;
memory[1628] <= 32'h0;
memory[1629] <= 32'h0;
memory[1630] <= 32'h0;
memory[1631] <= 32'h0;
memory[1632] <= 32'h0;
memory[1633] <= 32'h0;
memory[1634] <= 32'h0;
memory[1635] <= 32'h0;
memory[1636] <= 32'h0;
memory[1637] <= 32'h0;
memory[1638] <= 32'h0;
memory[1639] <= 32'h0;
memory[1640] <= 32'h0;
memory[1641] <= 32'h0;
memory[1642] <= 32'h0;
memory[1643] <= 32'h0;
memory[1644] <= 32'h0;
memory[1645] <= 32'h0;
memory[1646] <= 32'h0;
memory[1647] <= 32'h0;
memory[1648] <= 32'h0;
memory[1649] <= 32'h0;
memory[1650] <= 32'h0;
memory[1651] <= 32'h0;
memory[1652] <= 32'h0;
memory[1653] <= 32'h0;
memory[1654] <= 32'h0;
memory[1655] <= 32'h0;
memory[1656] <= 32'h0;
memory[1657] <= 32'h0;
memory[1658] <= 32'h0;
memory[1659] <= 32'h0;
memory[1660] <= 32'h0;
memory[1661] <= 32'h0;
memory[1662] <= 32'h0;
memory[1663] <= 32'h0;
memory[1664] <= 32'h0;
memory[1665] <= 32'h0;
memory[1666] <= 32'h0;
memory[1667] <= 32'h0;
memory[1668] <= 32'h0;
memory[1669] <= 32'h0;
memory[1670] <= 32'h0;
memory[1671] <= 32'h0;
memory[1672] <= 32'h0;
memory[1673] <= 32'h0;
memory[1674] <= 32'h0;
memory[1675] <= 32'h0;
memory[1676] <= 32'h0;
memory[1677] <= 32'h0;
memory[1678] <= 32'h0;
memory[1679] <= 32'h0;
memory[1680] <= 32'h0;
memory[1681] <= 32'h0;
memory[1682] <= 32'h0;
memory[1683] <= 32'h0;
memory[1684] <= 32'h0;
memory[1685] <= 32'h0;
memory[1686] <= 32'h0;
memory[1687] <= 32'h0;
memory[1688] <= 32'h0;
memory[1689] <= 32'h0;
memory[1690] <= 32'h0;
memory[1691] <= 32'h0;
memory[1692] <= 32'h0;
memory[1693] <= 32'h0;
memory[1694] <= 32'h0;
memory[1695] <= 32'h0;
memory[1696] <= 32'h0;
memory[1697] <= 32'h0;
memory[1698] <= 32'h0;
memory[1699] <= 32'h0;
memory[1700] <= 32'h0;
memory[1701] <= 32'h0;
memory[1702] <= 32'h0;
memory[1703] <= 32'h0;
memory[1704] <= 32'h0;
memory[1705] <= 32'h0;
memory[1706] <= 32'h0;
memory[1707] <= 32'h0;
memory[1708] <= 32'h0;
memory[1709] <= 32'h0;
memory[1710] <= 32'h0;
memory[1711] <= 32'h0;
memory[1712] <= 32'h0;
memory[1713] <= 32'h0;
memory[1714] <= 32'h0;
memory[1715] <= 32'h0;
memory[1716] <= 32'h0;
memory[1717] <= 32'h0;
memory[1718] <= 32'h0;
memory[1719] <= 32'h0;
memory[1720] <= 32'h0;
memory[1721] <= 32'h0;
memory[1722] <= 32'h0;
memory[1723] <= 32'h0;
memory[1724] <= 32'h0;
memory[1725] <= 32'h0;
memory[1726] <= 32'h0;
memory[1727] <= 32'h0;
memory[1728] <= 32'h0;
memory[1729] <= 32'h0;
memory[1730] <= 32'h0;
memory[1731] <= 32'h0;
memory[1732] <= 32'h0;
memory[1733] <= 32'h0;
memory[1734] <= 32'h0;
memory[1735] <= 32'h0;
memory[1736] <= 32'h0;
memory[1737] <= 32'h0;
memory[1738] <= 32'h0;
memory[1739] <= 32'h0;
memory[1740] <= 32'h0;
memory[1741] <= 32'h0;
memory[1742] <= 32'h0;
memory[1743] <= 32'h0;
memory[1744] <= 32'h0;
memory[1745] <= 32'h0;
memory[1746] <= 32'h0;
memory[1747] <= 32'h0;
memory[1748] <= 32'h0;
memory[1749] <= 32'h0;
memory[1750] <= 32'h0;
memory[1751] <= 32'h0;
memory[1752] <= 32'h0;
memory[1753] <= 32'h0;
memory[1754] <= 32'h0;
memory[1755] <= 32'h0;
memory[1756] <= 32'h0;
memory[1757] <= 32'h0;
memory[1758] <= 32'h0;
memory[1759] <= 32'h0;
memory[1760] <= 32'h0;
memory[1761] <= 32'h0;
memory[1762] <= 32'h0;
memory[1763] <= 32'h0;
memory[1764] <= 32'h0;
memory[1765] <= 32'h0;
memory[1766] <= 32'h0;
memory[1767] <= 32'h0;
memory[1768] <= 32'h0;
memory[1769] <= 32'h0;
memory[1770] <= 32'h0;
memory[1771] <= 32'h0;
memory[1772] <= 32'h0;
memory[1773] <= 32'h0;
memory[1774] <= 32'h0;
memory[1775] <= 32'h0;
memory[1776] <= 32'h0;
memory[1777] <= 32'h0;
memory[1778] <= 32'h0;
memory[1779] <= 32'h0;
memory[1780] <= 32'h0;
memory[1781] <= 32'h0;
memory[1782] <= 32'h0;
memory[1783] <= 32'h0;
memory[1784] <= 32'h0;
memory[1785] <= 32'h0;
memory[1786] <= 32'h0;
memory[1787] <= 32'h0;
memory[1788] <= 32'h0;
memory[1789] <= 32'h0;
memory[1790] <= 32'h0;
memory[1791] <= 32'h0;
memory[1792] <= 32'h0;
memory[1793] <= 32'h0;
memory[1794] <= 32'h0;
memory[1795] <= 32'h0;
memory[1796] <= 32'h0;
memory[1797] <= 32'h0;
memory[1798] <= 32'h0;
memory[1799] <= 32'h0;
memory[1800] <= 32'h0;
memory[1801] <= 32'h0;
memory[1802] <= 32'h0;
memory[1803] <= 32'h0;
memory[1804] <= 32'h0;
memory[1805] <= 32'h0;
memory[1806] <= 32'h0;
memory[1807] <= 32'h0;
memory[1808] <= 32'h0;
memory[1809] <= 32'h0;
memory[1810] <= 32'h0;
memory[1811] <= 32'h0;
memory[1812] <= 32'h0;
memory[1813] <= 32'h0;
memory[1814] <= 32'h0;
memory[1815] <= 32'h0;
memory[1816] <= 32'h0;
memory[1817] <= 32'h0;
memory[1818] <= 32'h0;
memory[1819] <= 32'h0;
memory[1820] <= 32'h0;
memory[1821] <= 32'h0;
memory[1822] <= 32'h0;
memory[1823] <= 32'h0;
memory[1824] <= 32'h0;
memory[1825] <= 32'h0;
memory[1826] <= 32'h0;
memory[1827] <= 32'h0;
memory[1828] <= 32'h0;
memory[1829] <= 32'h0;
memory[1830] <= 32'h0;
memory[1831] <= 32'h0;
memory[1832] <= 32'h0;
memory[1833] <= 32'h0;
memory[1834] <= 32'h0;
memory[1835] <= 32'h0;
memory[1836] <= 32'h0;
memory[1837] <= 32'h0;
memory[1838] <= 32'h0;
memory[1839] <= 32'h0;
memory[1840] <= 32'h0;
memory[1841] <= 32'h0;
memory[1842] <= 32'h0;
memory[1843] <= 32'h0;
memory[1844] <= 32'h0;
memory[1845] <= 32'h0;
memory[1846] <= 32'h0;
memory[1847] <= 32'h0;
memory[1848] <= 32'h0;
memory[1849] <= 32'h0;
memory[1850] <= 32'h0;
memory[1851] <= 32'h0;
memory[1852] <= 32'h0;
memory[1853] <= 32'h0;
memory[1854] <= 32'h0;
memory[1855] <= 32'h0;
memory[1856] <= 32'h0;
memory[1857] <= 32'h0;
memory[1858] <= 32'h0;
memory[1859] <= 32'h0;
memory[1860] <= 32'h0;
memory[1861] <= 32'h0;
memory[1862] <= 32'h0;
memory[1863] <= 32'h0;
memory[1864] <= 32'h0;
memory[1865] <= 32'h0;
memory[1866] <= 32'h0;
memory[1867] <= 32'h0;
memory[1868] <= 32'h0;
memory[1869] <= 32'h0;
memory[1870] <= 32'h0;
memory[1871] <= 32'h0;
memory[1872] <= 32'h0;
memory[1873] <= 32'h0;
memory[1874] <= 32'h0;
memory[1875] <= 32'h0;
memory[1876] <= 32'h0;
memory[1877] <= 32'h0;
memory[1878] <= 32'h0;
memory[1879] <= 32'h0;
memory[1880] <= 32'h0;
memory[1881] <= 32'h0;
memory[1882] <= 32'h0;
memory[1883] <= 32'h0;
memory[1884] <= 32'h0;
memory[1885] <= 32'h0;
memory[1886] <= 32'h0;
memory[1887] <= 32'h0;
memory[1888] <= 32'h0;
memory[1889] <= 32'h0;
memory[1890] <= 32'h0;
memory[1891] <= 32'h0;
memory[1892] <= 32'h0;
memory[1893] <= 32'h0;
memory[1894] <= 32'h0;
memory[1895] <= 32'h0;
memory[1896] <= 32'h0;
memory[1897] <= 32'h0;
memory[1898] <= 32'h0;
memory[1899] <= 32'h0;
memory[1900] <= 32'h0;
memory[1901] <= 32'h0;
memory[1902] <= 32'h0;
memory[1903] <= 32'h0;
memory[1904] <= 32'h0;
memory[1905] <= 32'h0;
memory[1906] <= 32'h0;
memory[1907] <= 32'h0;
memory[1908] <= 32'h0;
memory[1909] <= 32'h0;
memory[1910] <= 32'h0;
memory[1911] <= 32'h0;
memory[1912] <= 32'h0;
memory[1913] <= 32'h0;
memory[1914] <= 32'h0;
memory[1915] <= 32'h0;
memory[1916] <= 32'h0;
memory[1917] <= 32'h0;
memory[1918] <= 32'h0;
memory[1919] <= 32'h0;
memory[1920] <= 32'h0;
memory[1921] <= 32'h0;
memory[1922] <= 32'h0;
memory[1923] <= 32'h0;
memory[1924] <= 32'h0;
memory[1925] <= 32'h0;
memory[1926] <= 32'h0;
memory[1927] <= 32'h0;
memory[1928] <= 32'h0;
memory[1929] <= 32'h0;
memory[1930] <= 32'h0;
memory[1931] <= 32'h0;
memory[1932] <= 32'h0;
memory[1933] <= 32'h0;
memory[1934] <= 32'h0;
memory[1935] <= 32'h0;
memory[1936] <= 32'h0;
memory[1937] <= 32'h0;
memory[1938] <= 32'h0;
memory[1939] <= 32'h0;
memory[1940] <= 32'h0;
memory[1941] <= 32'h0;
memory[1942] <= 32'h0;
memory[1943] <= 32'h0;
memory[1944] <= 32'h0;
memory[1945] <= 32'h0;
memory[1946] <= 32'h0;
memory[1947] <= 32'h0;
memory[1948] <= 32'h0;
memory[1949] <= 32'h0;
memory[1950] <= 32'h0;
memory[1951] <= 32'h0;
memory[1952] <= 32'h0;
memory[1953] <= 32'h0;
memory[1954] <= 32'h0;
memory[1955] <= 32'h0;
memory[1956] <= 32'h0;
memory[1957] <= 32'h0;
memory[1958] <= 32'h0;
memory[1959] <= 32'h0;
memory[1960] <= 32'h0;
memory[1961] <= 32'h0;
memory[1962] <= 32'h0;
memory[1963] <= 32'h0;
memory[1964] <= 32'h0;
memory[1965] <= 32'h0;
memory[1966] <= 32'h0;
memory[1967] <= 32'h0;
memory[1968] <= 32'h0;
memory[1969] <= 32'h0;
memory[1970] <= 32'h0;
memory[1971] <= 32'h0;
memory[1972] <= 32'h0;
memory[1973] <= 32'h0;
memory[1974] <= 32'h0;
memory[1975] <= 32'h0;
memory[1976] <= 32'h0;
memory[1977] <= 32'h0;
memory[1978] <= 32'h0;
memory[1979] <= 32'h0;
memory[1980] <= 32'h0;
memory[1981] <= 32'h0;
memory[1982] <= 32'h0;
memory[1983] <= 32'h0;
memory[1984] <= 32'h0;
memory[1985] <= 32'h0;
memory[1986] <= 32'h0;
memory[1987] <= 32'h0;
memory[1988] <= 32'h0;
memory[1989] <= 32'h0;
memory[1990] <= 32'h0;
memory[1991] <= 32'h0;
memory[1992] <= 32'h0;
memory[1993] <= 32'h0;
memory[1994] <= 32'h0;
memory[1995] <= 32'h0;
memory[1996] <= 32'h0;
memory[1997] <= 32'h0;
memory[1998] <= 32'h0;
memory[1999] <= 32'h0;
memory[2000] <= 32'h0;
memory[2001] <= 32'h0;
memory[2002] <= 32'h0;
memory[2003] <= 32'h0;
memory[2004] <= 32'h0;
memory[2005] <= 32'h0;
memory[2006] <= 32'h0;
memory[2007] <= 32'h0;
memory[2008] <= 32'h0;
memory[2009] <= 32'h0;
memory[2010] <= 32'h0;
memory[2011] <= 32'h0;
memory[2012] <= 32'h0;
memory[2013] <= 32'h0;
memory[2014] <= 32'h0;
memory[2015] <= 32'h0;
memory[2016] <= 32'h0;
memory[2017] <= 32'h0;
memory[2018] <= 32'h0;
memory[2019] <= 32'h0;
memory[2020] <= 32'h0;
memory[2021] <= 32'h0;
memory[2022] <= 32'h0;
memory[2023] <= 32'h0;
memory[2024] <= 32'h0;
memory[2025] <= 32'h0;
memory[2026] <= 32'h0;
memory[2027] <= 32'h0;
memory[2028] <= 32'h0;
memory[2029] <= 32'h0;
memory[2030] <= 32'h0;
memory[2031] <= 32'h0;
memory[2032] <= 32'h0;
memory[2033] <= 32'h0;
memory[2034] <= 32'h0;
memory[2035] <= 32'h0;
memory[2036] <= 32'h0;
memory[2037] <= 32'h0;
memory[2038] <= 32'h0;
memory[2039] <= 32'h0;
memory[2040] <= 32'h0;
memory[2041] <= 32'h0;
memory[2042] <= 32'h0;
memory[2043] <= 32'h0;
memory[2044] <= 32'h0;
memory[2045] <= 32'h0;
memory[2046] <= 32'h0;
memory[2047] <= 32'h0;
memory[2048] <= 32'h0;
memory[2049] <= 32'h0;
memory[2050] <= 32'h0;
memory[2051] <= 32'h0;
memory[2052] <= 32'h0;
memory[2053] <= 32'h0;
memory[2054] <= 32'h0;
memory[2055] <= 32'h0;
memory[2056] <= 32'h0;
memory[2057] <= 32'h0;
memory[2058] <= 32'h0;
memory[2059] <= 32'h0;
memory[2060] <= 32'h0;
memory[2061] <= 32'h0;
memory[2062] <= 32'h0;
memory[2063] <= 32'h0;
memory[2064] <= 32'h0;
memory[2065] <= 32'h0;
memory[2066] <= 32'h0;
memory[2067] <= 32'h0;
memory[2068] <= 32'h0;
memory[2069] <= 32'h0;
memory[2070] <= 32'h0;
memory[2071] <= 32'h0;
memory[2072] <= 32'h0;
memory[2073] <= 32'h0;
memory[2074] <= 32'h0;
memory[2075] <= 32'h0;
memory[2076] <= 32'h0;
memory[2077] <= 32'h0;
memory[2078] <= 32'h0;
memory[2079] <= 32'h0;
memory[2080] <= 32'h0;
memory[2081] <= 32'h0;
memory[2082] <= 32'h0;
memory[2083] <= 32'h0;
memory[2084] <= 32'h0;
memory[2085] <= 32'h0;
memory[2086] <= 32'h0;
memory[2087] <= 32'h0;
memory[2088] <= 32'h0;
memory[2089] <= 32'h0;
memory[2090] <= 32'h0;
memory[2091] <= 32'h0;
memory[2092] <= 32'h0;
memory[2093] <= 32'h0;
memory[2094] <= 32'h0;
memory[2095] <= 32'h0;
memory[2096] <= 32'h0;
memory[2097] <= 32'h0;
memory[2098] <= 32'h0;
memory[2099] <= 32'h0;
memory[2100] <= 32'h0;
memory[2101] <= 32'h0;
memory[2102] <= 32'h0;
memory[2103] <= 32'h0;
memory[2104] <= 32'h0;
memory[2105] <= 32'h0;
memory[2106] <= 32'h0;
memory[2107] <= 32'h0;
memory[2108] <= 32'h0;
memory[2109] <= 32'h0;
memory[2110] <= 32'h0;
memory[2111] <= 32'h0;
memory[2112] <= 32'h0;
memory[2113] <= 32'h0;
memory[2114] <= 32'h0;
memory[2115] <= 32'h0;
memory[2116] <= 32'h0;
memory[2117] <= 32'h0;
memory[2118] <= 32'h0;
memory[2119] <= 32'h0;
memory[2120] <= 32'h0;
memory[2121] <= 32'h0;
memory[2122] <= 32'h0;
memory[2123] <= 32'h0;
memory[2124] <= 32'h0;
memory[2125] <= 32'h0;
memory[2126] <= 32'h0;
memory[2127] <= 32'h0;
memory[2128] <= 32'h0;
memory[2129] <= 32'h0;
memory[2130] <= 32'h0;
memory[2131] <= 32'h0;
memory[2132] <= 32'h0;
memory[2133] <= 32'h0;
memory[2134] <= 32'h0;
memory[2135] <= 32'h0;
memory[2136] <= 32'h0;
memory[2137] <= 32'h0;
memory[2138] <= 32'h0;
memory[2139] <= 32'h0;
memory[2140] <= 32'h0;
memory[2141] <= 32'h0;
memory[2142] <= 32'h0;
memory[2143] <= 32'h0;
memory[2144] <= 32'h0;
memory[2145] <= 32'h0;
memory[2146] <= 32'h0;
memory[2147] <= 32'h0;
memory[2148] <= 32'h0;
memory[2149] <= 32'h0;
memory[2150] <= 32'h0;
memory[2151] <= 32'h0;
memory[2152] <= 32'h0;
memory[2153] <= 32'h0;
memory[2154] <= 32'h0;
memory[2155] <= 32'h0;
memory[2156] <= 32'h0;
memory[2157] <= 32'h0;
memory[2158] <= 32'h0;
memory[2159] <= 32'h0;
memory[2160] <= 32'h0;
memory[2161] <= 32'h0;
memory[2162] <= 32'h0;
memory[2163] <= 32'h0;
memory[2164] <= 32'h0;
memory[2165] <= 32'h0;
memory[2166] <= 32'h0;
memory[2167] <= 32'h0;
memory[2168] <= 32'h0;
memory[2169] <= 32'h0;
memory[2170] <= 32'h0;
memory[2171] <= 32'h0;
memory[2172] <= 32'h0;
memory[2173] <= 32'h0;
memory[2174] <= 32'h0;
memory[2175] <= 32'h0;
memory[2176] <= 32'h0;
memory[2177] <= 32'h0;
memory[2178] <= 32'h0;
memory[2179] <= 32'h0;
memory[2180] <= 32'h0;
memory[2181] <= 32'h0;
memory[2182] <= 32'h0;
memory[2183] <= 32'h0;
memory[2184] <= 32'h0;
memory[2185] <= 32'h0;
memory[2186] <= 32'h0;
memory[2187] <= 32'h0;
memory[2188] <= 32'h0;
memory[2189] <= 32'h0;
memory[2190] <= 32'h0;
memory[2191] <= 32'h0;
memory[2192] <= 32'h0;
memory[2193] <= 32'h0;
memory[2194] <= 32'h0;
memory[2195] <= 32'h0;
memory[2196] <= 32'h0;
memory[2197] <= 32'h0;
memory[2198] <= 32'h0;
memory[2199] <= 32'h0;
memory[2200] <= 32'h0;
memory[2201] <= 32'h0;
memory[2202] <= 32'h0;
memory[2203] <= 32'h0;
memory[2204] <= 32'h0;
memory[2205] <= 32'h0;
memory[2206] <= 32'h0;
memory[2207] <= 32'h0;
memory[2208] <= 32'h0;
memory[2209] <= 32'h0;
memory[2210] <= 32'h0;
memory[2211] <= 32'h0;
memory[2212] <= 32'h0;
memory[2213] <= 32'h0;
memory[2214] <= 32'h0;
memory[2215] <= 32'h0;
memory[2216] <= 32'h0;
memory[2217] <= 32'h0;
memory[2218] <= 32'h0;
memory[2219] <= 32'h0;
memory[2220] <= 32'h0;
memory[2221] <= 32'h0;
memory[2222] <= 32'h0;
memory[2223] <= 32'h0;
memory[2224] <= 32'h0;
memory[2225] <= 32'h0;
memory[2226] <= 32'h0;
memory[2227] <= 32'h0;
memory[2228] <= 32'h0;
memory[2229] <= 32'h0;
memory[2230] <= 32'h0;
memory[2231] <= 32'h0;
memory[2232] <= 32'h0;
memory[2233] <= 32'h0;
memory[2234] <= 32'h0;
memory[2235] <= 32'h0;
memory[2236] <= 32'h0;
memory[2237] <= 32'h0;
memory[2238] <= 32'h0;
memory[2239] <= 32'h0;
memory[2240] <= 32'h0;
memory[2241] <= 32'h0;
memory[2242] <= 32'h0;
memory[2243] <= 32'h0;
memory[2244] <= 32'h0;
memory[2245] <= 32'h0;
memory[2246] <= 32'h0;
memory[2247] <= 32'h0;
memory[2248] <= 32'h0;
memory[2249] <= 32'h0;
memory[2250] <= 32'h0;
memory[2251] <= 32'h0;
memory[2252] <= 32'h0;
memory[2253] <= 32'h0;
memory[2254] <= 32'h0;
memory[2255] <= 32'h0;
memory[2256] <= 32'h0;
memory[2257] <= 32'h0;
memory[2258] <= 32'h0;
memory[2259] <= 32'h0;
memory[2260] <= 32'h0;
memory[2261] <= 32'h0;
memory[2262] <= 32'h0;
memory[2263] <= 32'h0;
memory[2264] <= 32'h0;
memory[2265] <= 32'h0;
memory[2266] <= 32'h0;
memory[2267] <= 32'h0;
memory[2268] <= 32'h0;
memory[2269] <= 32'h0;
memory[2270] <= 32'h0;
memory[2271] <= 32'h0;
memory[2272] <= 32'h0;
memory[2273] <= 32'h0;
memory[2274] <= 32'h0;
memory[2275] <= 32'h0;
memory[2276] <= 32'h0;
memory[2277] <= 32'h0;
memory[2278] <= 32'h0;
memory[2279] <= 32'h0;
memory[2280] <= 32'h0;
memory[2281] <= 32'h0;
memory[2282] <= 32'h0;
memory[2283] <= 32'h0;
memory[2284] <= 32'h0;
memory[2285] <= 32'h0;
memory[2286] <= 32'h0;
memory[2287] <= 32'h0;
memory[2288] <= 32'h0;
memory[2289] <= 32'h0;
memory[2290] <= 32'h0;
memory[2291] <= 32'h0;
memory[2292] <= 32'h0;
memory[2293] <= 32'h0;
memory[2294] <= 32'h0;
memory[2295] <= 32'h0;
memory[2296] <= 32'h0;
memory[2297] <= 32'h0;
memory[2298] <= 32'h0;
memory[2299] <= 32'h0;
memory[2300] <= 32'h0;
memory[2301] <= 32'h0;
memory[2302] <= 32'h0;
memory[2303] <= 32'h0;
memory[2304] <= 32'h0;
memory[2305] <= 32'h0;
memory[2306] <= 32'h0;
memory[2307] <= 32'h0;
memory[2308] <= 32'h0;
memory[2309] <= 32'h0;
memory[2310] <= 32'h0;
memory[2311] <= 32'h0;
memory[2312] <= 32'h0;
memory[2313] <= 32'h0;
memory[2314] <= 32'h0;
memory[2315] <= 32'h0;
memory[2316] <= 32'h0;
memory[2317] <= 32'h0;
memory[2318] <= 32'h0;
memory[2319] <= 32'h0;
memory[2320] <= 32'h0;
memory[2321] <= 32'h0;
memory[2322] <= 32'h0;
memory[2323] <= 32'h0;
memory[2324] <= 32'h0;
memory[2325] <= 32'h0;
memory[2326] <= 32'h0;
memory[2327] <= 32'h0;
memory[2328] <= 32'h0;
memory[2329] <= 32'h0;
memory[2330] <= 32'h0;
memory[2331] <= 32'h0;
memory[2332] <= 32'h0;
memory[2333] <= 32'h0;
memory[2334] <= 32'h0;
memory[2335] <= 32'h0;
memory[2336] <= 32'h0;
memory[2337] <= 32'h0;
memory[2338] <= 32'h0;
memory[2339] <= 32'h0;
memory[2340] <= 32'h0;
memory[2341] <= 32'h0;
memory[2342] <= 32'h0;
memory[2343] <= 32'h0;
memory[2344] <= 32'h0;
memory[2345] <= 32'h0;
memory[2346] <= 32'h0;
memory[2347] <= 32'h0;
memory[2348] <= 32'h0;
memory[2349] <= 32'h0;
memory[2350] <= 32'h0;
memory[2351] <= 32'h0;
memory[2352] <= 32'h0;
memory[2353] <= 32'h0;
memory[2354] <= 32'h0;
memory[2355] <= 32'h0;
memory[2356] <= 32'h0;
memory[2357] <= 32'h0;
memory[2358] <= 32'h0;
memory[2359] <= 32'h0;
memory[2360] <= 32'h0;
memory[2361] <= 32'h0;
memory[2362] <= 32'h0;
memory[2363] <= 32'h0;
memory[2364] <= 32'h0;
memory[2365] <= 32'h0;
memory[2366] <= 32'h0;
memory[2367] <= 32'h0;
memory[2368] <= 32'h0;
memory[2369] <= 32'h0;
memory[2370] <= 32'h0;
memory[2371] <= 32'h0;
memory[2372] <= 32'h0;
memory[2373] <= 32'h0;
memory[2374] <= 32'h0;
memory[2375] <= 32'h0;
memory[2376] <= 32'h0;
memory[2377] <= 32'h0;
memory[2378] <= 32'h0;
memory[2379] <= 32'h0;
memory[2380] <= 32'h0;
memory[2381] <= 32'h0;
memory[2382] <= 32'h0;
memory[2383] <= 32'h0;
memory[2384] <= 32'h0;
memory[2385] <= 32'h0;
memory[2386] <= 32'h0;
memory[2387] <= 32'h0;
memory[2388] <= 32'h0;
memory[2389] <= 32'h0;
memory[2390] <= 32'h0;
memory[2391] <= 32'h0;
memory[2392] <= 32'h0;
memory[2393] <= 32'h0;
memory[2394] <= 32'h0;
memory[2395] <= 32'h0;
memory[2396] <= 32'h0;
memory[2397] <= 32'h0;
memory[2398] <= 32'h0;
memory[2399] <= 32'h0;
memory[2400] <= 32'h0;
memory[2401] <= 32'h0;
memory[2402] <= 32'h0;
memory[2403] <= 32'h0;
memory[2404] <= 32'h0;
memory[2405] <= 32'h0;
memory[2406] <= 32'h0;
memory[2407] <= 32'h0;
memory[2408] <= 32'h0;
memory[2409] <= 32'h0;
memory[2410] <= 32'h0;
memory[2411] <= 32'h0;
memory[2412] <= 32'h0;
memory[2413] <= 32'h0;
memory[2414] <= 32'h0;
memory[2415] <= 32'h0;
memory[2416] <= 32'h0;
memory[2417] <= 32'h0;
memory[2418] <= 32'h0;
memory[2419] <= 32'h0;
memory[2420] <= 32'h0;
memory[2421] <= 32'h0;
memory[2422] <= 32'h0;
memory[2423] <= 32'h0;
memory[2424] <= 32'h0;
memory[2425] <= 32'h0;
memory[2426] <= 32'h0;
memory[2427] <= 32'h0;
memory[2428] <= 32'h0;
memory[2429] <= 32'h0;
memory[2430] <= 32'h0;
memory[2431] <= 32'h0;
memory[2432] <= 32'h0;
memory[2433] <= 32'h0;
memory[2434] <= 32'h0;
memory[2435] <= 32'h0;
memory[2436] <= 32'h0;
memory[2437] <= 32'h0;
memory[2438] <= 32'h0;
memory[2439] <= 32'h0;
memory[2440] <= 32'h0;
memory[2441] <= 32'h0;
memory[2442] <= 32'h0;
memory[2443] <= 32'h0;
memory[2444] <= 32'h0;
memory[2445] <= 32'h0;
memory[2446] <= 32'h0;
memory[2447] <= 32'h0;
memory[2448] <= 32'h0;
memory[2449] <= 32'h0;
memory[2450] <= 32'h0;
memory[2451] <= 32'h0;
memory[2452] <= 32'h0;
memory[2453] <= 32'h0;
memory[2454] <= 32'h0;
memory[2455] <= 32'h0;
memory[2456] <= 32'h0;
memory[2457] <= 32'h0;
memory[2458] <= 32'h0;
memory[2459] <= 32'h0;
memory[2460] <= 32'h0;
memory[2461] <= 32'h0;
memory[2462] <= 32'h0;
memory[2463] <= 32'h0;
memory[2464] <= 32'h0;
memory[2465] <= 32'h0;
memory[2466] <= 32'h0;
memory[2467] <= 32'h0;
memory[2468] <= 32'h0;
memory[2469] <= 32'h0;
memory[2470] <= 32'h0;
memory[2471] <= 32'h0;
memory[2472] <= 32'h0;
memory[2473] <= 32'h0;
memory[2474] <= 32'h0;
memory[2475] <= 32'h0;
memory[2476] <= 32'h0;
memory[2477] <= 32'h0;
memory[2478] <= 32'h0;
memory[2479] <= 32'h0;
memory[2480] <= 32'h0;
memory[2481] <= 32'h0;
memory[2482] <= 32'h0;
memory[2483] <= 32'h0;
memory[2484] <= 32'h0;
memory[2485] <= 32'h0;
memory[2486] <= 32'h0;
memory[2487] <= 32'h0;
memory[2488] <= 32'h0;
memory[2489] <= 32'h0;
memory[2490] <= 32'h0;
memory[2491] <= 32'h0;
memory[2492] <= 32'h0;
memory[2493] <= 32'h0;
memory[2494] <= 32'h0;
memory[2495] <= 32'h0;
memory[2496] <= 32'h0;
memory[2497] <= 32'h0;
memory[2498] <= 32'h0;
memory[2499] <= 32'h0;
memory[2500] <= 32'h0;
memory[2501] <= 32'h0;
memory[2502] <= 32'h0;
memory[2503] <= 32'h0;
memory[2504] <= 32'h0;
memory[2505] <= 32'h0;
memory[2506] <= 32'h0;
memory[2507] <= 32'h0;
memory[2508] <= 32'h0;
memory[2509] <= 32'h0;
memory[2510] <= 32'h0;
memory[2511] <= 32'h0;
memory[2512] <= 32'h0;
memory[2513] <= 32'h0;
memory[2514] <= 32'h0;
memory[2515] <= 32'h0;
memory[2516] <= 32'h0;
memory[2517] <= 32'h0;
memory[2518] <= 32'h0;
memory[2519] <= 32'h0;
memory[2520] <= 32'h0;
memory[2521] <= 32'h0;
memory[2522] <= 32'h0;
memory[2523] <= 32'h0;
memory[2524] <= 32'h0;
memory[2525] <= 32'h0;
memory[2526] <= 32'h0;
memory[2527] <= 32'h0;
memory[2528] <= 32'h0;
memory[2529] <= 32'h0;
memory[2530] <= 32'h0;
memory[2531] <= 32'h0;
memory[2532] <= 32'h0;
memory[2533] <= 32'h0;
memory[2534] <= 32'h0;
memory[2535] <= 32'h0;
memory[2536] <= 32'h0;
memory[2537] <= 32'h0;
memory[2538] <= 32'h0;
memory[2539] <= 32'h0;
memory[2540] <= 32'h0;
memory[2541] <= 32'h0;
memory[2542] <= 32'h0;
memory[2543] <= 32'h0;
memory[2544] <= 32'h0;
memory[2545] <= 32'h0;
memory[2546] <= 32'h0;
memory[2547] <= 32'h0;
memory[2548] <= 32'h0;
memory[2549] <= 32'h0;
memory[2550] <= 32'h0;
memory[2551] <= 32'h1;
memory[2552] <= 32'h1;
memory[2553] <= 32'h1;
memory[2554] <= 32'h1;
memory[2555] <= 32'h0;
memory[2556] <= 32'h0;
memory[2557] <= 32'h0;
memory[2558] <= 32'h0;
memory[2559] <= 32'h0;
memory[2560] <= 32'h0;
memory[2561] <= 32'h0;
memory[2562] <= 32'h0;
memory[2563] <= 32'h0;
memory[2564] <= 32'h0;
memory[2565] <= 32'h0;
memory[2566] <= 32'h0;
memory[2567] <= 32'h0;
memory[2568] <= 32'h0;
memory[2569] <= 32'h0;
memory[2570] <= 32'h0;
memory[2571] <= 32'h0;
memory[2572] <= 32'h0;
memory[2573] <= 32'h0;
memory[2574] <= 32'h0;
memory[2575] <= 32'h0;
memory[2576] <= 32'h0;
memory[2577] <= 32'h0;
memory[2578] <= 32'h0;
memory[2579] <= 32'h0;
memory[2580] <= 32'h0;
memory[2581] <= 32'h0;
memory[2582] <= 32'h1;
memory[2583] <= 32'h1;
memory[2584] <= 32'h1;
memory[2585] <= 32'h1;
memory[2586] <= 32'h0;
memory[2587] <= 32'h0;
memory[2588] <= 32'h0;
memory[2589] <= 32'h0;
memory[2590] <= 32'h0;
memory[2591] <= 32'h0;
memory[2592] <= 32'h0;
memory[2593] <= 32'h0;
memory[2594] <= 32'h0;
memory[2595] <= 32'h0;
memory[2596] <= 32'h0;
memory[2597] <= 32'h0;
memory[2598] <= 32'h0;
memory[2599] <= 32'h0;
memory[2600] <= 32'h0;
memory[2601] <= 32'h0;
memory[2602] <= 32'h0;
memory[2603] <= 32'h0;
memory[2604] <= 32'h0;
memory[2605] <= 32'h0;
memory[2606] <= 32'h0;
memory[2607] <= 32'h0;
memory[2608] <= 32'h0;
memory[2609] <= 32'h0;
memory[2610] <= 32'h0;
memory[2611] <= 32'h0;
memory[2612] <= 32'h0;
memory[2613] <= 32'h1;
memory[2614] <= 32'h1;
memory[2615] <= 32'h1;
memory[2616] <= 32'h1;
memory[2617] <= 32'h0;
memory[2618] <= 32'h0;
memory[2619] <= 32'h0;
memory[2620] <= 32'h0;
memory[2621] <= 32'h0;
memory[2622] <= 32'h0;
memory[2623] <= 32'h0;
memory[2624] <= 32'h0;
memory[2625] <= 32'h0;
memory[2626] <= 32'h0;
memory[2627] <= 32'h0;
memory[2628] <= 32'h0;
memory[2629] <= 32'h0;
memory[2630] <= 32'h0;
memory[2631] <= 32'h0;
memory[2632] <= 32'h0;
memory[2633] <= 32'h0;
memory[2634] <= 32'h0;
memory[2635] <= 32'h0;
memory[2636] <= 32'h0;
memory[2637] <= 32'h0;
memory[2638] <= 32'h0;
memory[2639] <= 32'h0;
memory[2640] <= 32'h0;
memory[2641] <= 32'h0;
memory[2642] <= 32'h0;
memory[2643] <= 32'h0;
memory[2644] <= 32'h1;
memory[2645] <= 32'h1;
memory[2646] <= 32'h1;
memory[2647] <= 32'h1;
memory[2648] <= 32'h0;
memory[2649] <= 32'h0;
memory[2650] <= 32'h0;
memory[2651] <= 32'h0;
memory[2652] <= 32'h0;
memory[2653] <= 32'h0;
memory[2654] <= 32'h0;
memory[2655] <= 32'h0;
memory[2656] <= 32'h0;
memory[2657] <= 32'h0;
memory[2658] <= 32'h0;
memory[2659] <= 32'h0;
memory[2660] <= 32'h0;
memory[2661] <= 32'h0;
memory[2662] <= 32'h0;
memory[2663] <= 32'h0;
memory[2664] <= 32'h0;
memory[2665] <= 32'h0;
memory[2666] <= 32'h0;
memory[2667] <= 32'h0;
memory[2668] <= 32'h0;
memory[2669] <= 32'h0;
memory[2670] <= 32'h0;
memory[2671] <= 32'h0;
memory[2672] <= 32'h0;
memory[2673] <= 32'h0;
memory[2674] <= 32'h0;
memory[2675] <= 32'h1;
memory[2676] <= 32'h1;
memory[2677] <= 32'h1;
memory[2678] <= 32'h1;
memory[2679] <= 32'h0;
memory[2680] <= 32'h0;
memory[2681] <= 32'h0;
memory[2682] <= 32'h0;
memory[2683] <= 32'h0;
memory[2684] <= 32'h0;
memory[2685] <= 32'h0;
memory[2686] <= 32'h0;
memory[2687] <= 32'h0;
memory[2688] <= 32'h0;
memory[2689] <= 32'h0;
memory[2690] <= 32'h0;
memory[2691] <= 32'h0;
memory[2692] <= 32'h0;
memory[2693] <= 32'h0;
memory[2694] <= 32'h0;
memory[2695] <= 32'h0;
memory[2696] <= 32'h0;
memory[2697] <= 32'h0;
memory[2698] <= 32'h0;
memory[2699] <= 32'h0;
memory[2700] <= 32'h0;
memory[2701] <= 32'h0;
memory[2702] <= 32'h0;
memory[2703] <= 32'h0;
memory[2704] <= 32'h0;
memory[2705] <= 32'h0;
memory[2706] <= 32'h1;
memory[2707] <= 32'h1;
memory[2708] <= 32'h1;
memory[2709] <= 32'h1;
memory[2710] <= 32'h0;
memory[2711] <= 32'h0;
memory[2712] <= 32'h0;
memory[2713] <= 32'h0;
memory[2714] <= 32'h0;
memory[2715] <= 32'h0;
memory[2716] <= 32'h0;
memory[2717] <= 32'h0;
memory[2718] <= 32'h0;
memory[2719] <= 32'h0;
memory[2720] <= 32'h0;
memory[2721] <= 32'h0;
memory[2722] <= 32'h0;
memory[2723] <= 32'h0;
memory[2724] <= 32'h0;
memory[2725] <= 32'h0;
memory[2726] <= 32'h0;
memory[2727] <= 32'h0;
memory[2728] <= 32'h0;
memory[2729] <= 32'h0;
memory[2730] <= 32'h0;
memory[2731] <= 32'h0;
memory[2732] <= 32'h0;
memory[2733] <= 32'h0;
memory[2734] <= 32'h0;
memory[2735] <= 32'h0;
memory[2736] <= 32'h0;
memory[2737] <= 32'h1;
memory[2738] <= 32'h1;
memory[2739] <= 32'h1;
memory[2740] <= 32'h1;
memory[2741] <= 32'h0;
memory[2742] <= 32'h0;
memory[2743] <= 32'h0;
memory[2744] <= 32'h0;
memory[2745] <= 32'h0;
memory[2746] <= 32'h0;
memory[2747] <= 32'h0;
memory[2748] <= 32'h0;
memory[2749] <= 32'h0;
memory[2750] <= 32'h0;
memory[2751] <= 32'h0;
memory[2752] <= 32'h0;
memory[2753] <= 32'h0;
memory[2754] <= 32'h0;
memory[2755] <= 32'h0;
memory[2756] <= 32'h0;
memory[2757] <= 32'h0;
memory[2758] <= 32'h0;
memory[2759] <= 32'h0;
memory[2760] <= 32'h0;
memory[2761] <= 32'h0;
memory[2762] <= 32'h0;
memory[2763] <= 32'h0;
memory[2764] <= 32'h0;
memory[2765] <= 32'h0;
memory[2766] <= 32'h0;
memory[2767] <= 32'h0;
memory[2768] <= 32'h1;
memory[2769] <= 32'h1;
memory[2770] <= 32'h1;
memory[2771] <= 32'h1;
memory[2772] <= 32'h0;
memory[2773] <= 32'h0;
memory[2774] <= 32'h0;
memory[2775] <= 32'h0;
memory[2776] <= 32'h0;
memory[2777] <= 32'h0;
memory[2778] <= 32'h0;
memory[2779] <= 32'h0;
memory[2780] <= 32'h0;
memory[2781] <= 32'h0;
memory[2782] <= 32'h0;
memory[2783] <= 32'h0;
memory[2784] <= 32'h0;
memory[2785] <= 32'h0;
memory[2786] <= 32'h0;
memory[2787] <= 32'h0;
memory[2788] <= 32'h0;
memory[2789] <= 32'h0;
memory[2790] <= 32'h0;
memory[2791] <= 32'h0;
memory[2792] <= 32'h0;
memory[2793] <= 32'h0;
memory[2794] <= 32'h0;
memory[2795] <= 32'h0;
memory[2796] <= 32'h0;
memory[2797] <= 32'h0;
memory[2798] <= 32'h0;
memory[2799] <= 32'h1;
memory[2800] <= 32'h1;
memory[2801] <= 32'h1;
memory[2802] <= 32'h1;
memory[2803] <= 32'h1;
memory[2804] <= 32'h1;
memory[2805] <= 32'h1;
memory[2806] <= 32'h1;
memory[2807] <= 32'h1;
memory[2808] <= 32'h1;
memory[2809] <= 32'h1;
memory[2810] <= 32'h1;
memory[2811] <= 32'h1;
memory[2812] <= 32'h1;
memory[2813] <= 32'h1;
memory[2814] <= 32'h1;
memory[2815] <= 32'h1;
memory[2816] <= 32'h1;
memory[2817] <= 32'h1;
memory[2818] <= 32'h1;
memory[2819] <= 32'h1;
memory[2820] <= 32'h1;
memory[2821] <= 32'h1;
memory[2822] <= 32'h1;
memory[2823] <= 32'h1;
memory[2824] <= 32'h1;
memory[2825] <= 32'h1;
memory[2826] <= 32'h1;
memory[2827] <= 32'h1;
memory[2828] <= 32'h1;
memory[2829] <= 32'h1;
memory[2830] <= 32'h1;
memory[2831] <= 32'h13;
memory[2832] <= 32'h20;
memory[2833] <= 32'h4;
memory[2834] <= 32'h4;
memory[2835] <= 32'h1;
memory[2836] <= 32'h1;
memory[2837] <= 32'h1;
memory[2838] <= 32'h1;
memory[2839] <= 32'h0;
memory[2840] <= 32'h0;
memory[2841] <= 32'h0;
memory[2842] <= 32'h0;
memory[2843] <= 32'h0;
memory[2844] <= 32'h0;
memory[2845] <= 32'h0;
memory[2846] <= 32'h0;
memory[2847] <= 32'h0;
memory[2848] <= 32'h0;
memory[2849] <= 32'h0;
memory[2850] <= 32'h0;
memory[2851] <= 32'h0;
memory[2852] <= 32'h0;
memory[2853] <= 32'h0;
memory[2854] <= 32'h0;
memory[2855] <= 32'h0;
memory[2856] <= 32'h0;
memory[2857] <= 32'h0;
memory[2858] <= 32'h0;
memory[2859] <= 32'h0;
memory[2860] <= 32'h0;
memory[2861] <= 32'h0;
memory[2862] <= 32'h0;
memory[2863] <= 32'h0;
memory[2864] <= 32'h0;
memory[2865] <= 32'h0;
memory[2866] <= 32'h0;
memory[2867] <= 32'h1;
memory[2868] <= 32'h1;
memory[2869] <= 32'h1;
memory[2870] <= 32'h1;
memory[2871] <= 32'h0;
memory[2872] <= 32'h0;
memory[2873] <= 32'h0;
memory[2874] <= 32'h0;
memory[2875] <= 32'h0;
memory[2876] <= 32'h0;
memory[2877] <= 32'h0;
memory[2878] <= 32'h0;
memory[2879] <= 32'h0;
memory[2880] <= 32'h0;
memory[2881] <= 32'h0;
memory[2882] <= 32'h0;
memory[2883] <= 32'h0;
memory[2884] <= 32'h0;
memory[2885] <= 32'h0;
memory[2886] <= 32'h0;
memory[2887] <= 32'h0;
memory[2888] <= 32'h0;
memory[2889] <= 32'h0;
memory[2890] <= 32'h0;
memory[2891] <= 32'h0;
memory[2892] <= 32'h0;
memory[2893] <= 32'h0;
memory[2894] <= 32'h0;
memory[2895] <= 32'h0;
memory[2896] <= 32'h0;
memory[2897] <= 32'h0;
memory[2898] <= 32'h0;
memory[2899] <= 32'h1;
memory[2900] <= 32'h1;
memory[2901] <= 32'h1;
memory[2902] <= 32'h1;
memory[2903] <= 32'h0;
memory[2904] <= 32'h0;
memory[2905] <= 32'h0;
memory[2906] <= 32'h0;
memory[2907] <= 32'h0;
memory[2908] <= 32'h0;
memory[2909] <= 32'h0;
memory[2910] <= 32'h0;
memory[2911] <= 32'h0;
memory[2912] <= 32'h0;
memory[2913] <= 32'h0;
memory[2914] <= 32'h0;
memory[2915] <= 32'h0;
memory[2916] <= 32'h0;
memory[2917] <= 32'h0;
memory[2918] <= 32'h0;
memory[2919] <= 32'h0;
memory[2920] <= 32'h0;
memory[2921] <= 32'h0;
memory[2922] <= 32'h0;
memory[2923] <= 32'h0;
memory[2924] <= 32'h0;
memory[2925] <= 32'h0;
memory[2926] <= 32'h0;
memory[2927] <= 32'h0;
memory[2928] <= 32'h0;
memory[2929] <= 32'h0;
memory[2930] <= 32'h0;
memory[2931] <= 32'h1;
memory[2932] <= 32'h1;
memory[2933] <= 32'h1;
memory[2934] <= 32'h1;
memory[2935] <= 32'h0;
memory[2936] <= 32'h0;
memory[2937] <= 32'h0;
memory[2938] <= 32'h0;
memory[2939] <= 32'h0;
memory[2940] <= 32'h0;
memory[2941] <= 32'h0;
memory[2942] <= 32'h0;
memory[2943] <= 32'h0;
memory[2944] <= 32'h0;
memory[2945] <= 32'h0;
memory[2946] <= 32'h0;
memory[2947] <= 32'h0;
memory[2948] <= 32'h0;
memory[2949] <= 32'h0;
memory[2950] <= 32'h0;
memory[2951] <= 32'h0;
memory[2952] <= 32'h0;
memory[2953] <= 32'h0;
memory[2954] <= 32'h0;
memory[2955] <= 32'h0;
memory[2956] <= 32'h0;
memory[2957] <= 32'h0;
memory[2958] <= 32'h0;
memory[2959] <= 32'h0;
memory[2960] <= 32'h0;
memory[2961] <= 32'h0;
memory[2962] <= 32'h0;
memory[2963] <= 32'h0;
memory[2964] <= 32'h0;
memory[2965] <= 32'h0;
memory[2966] <= 32'h0;
memory[2967] <= 32'h0;
memory[2968] <= 32'h0;
memory[2969] <= 32'h0;
memory[2970] <= 32'h0;
memory[2971] <= 32'h0;
memory[2972] <= 32'h0;
memory[2973] <= 32'h0;
memory[2974] <= 32'h0;
memory[2975] <= 32'h0;
memory[2976] <= 32'h0;
memory[2977] <= 32'h0;
memory[2978] <= 32'h0;
memory[2979] <= 32'h0;
memory[2980] <= 32'h0;
memory[2981] <= 32'h0;
memory[2982] <= 32'h0;
memory[2983] <= 32'h0;
memory[2984] <= 32'h0;
memory[2985] <= 32'h0;
memory[2986] <= 32'h0;
memory[2987] <= 32'h0;
memory[2988] <= 32'h0;
memory[2989] <= 32'h0;
memory[2990] <= 32'h0;
memory[2991] <= 32'h0;
memory[2992] <= 32'h0;
memory[2993] <= 32'h0;
memory[2994] <= 32'h0;
memory[2995] <= 32'h0;
memory[2996] <= 32'h0;
memory[2997] <= 32'h0;
memory[2998] <= 32'h0;
memory[2999] <= 32'h0;
memory[3000] <= 32'h0;
memory[3001] <= 32'h0;
memory[3002] <= 32'h0;
memory[3003] <= 32'h0;
memory[3004] <= 32'h0;
memory[3005] <= 32'h0;
memory[3006] <= 32'h0;
memory[3007] <= 32'h0;
memory[3008] <= 32'h0;
memory[3009] <= 32'h0;
memory[3010] <= 32'h0;
memory[3011] <= 32'h0;
memory[3012] <= 32'h0;
memory[3013] <= 32'h0;
memory[3014] <= 32'h0;
memory[3015] <= 32'h0;
memory[3016] <= 32'h0;
memory[3017] <= 32'h0;
memory[3018] <= 32'h0;
memory[3019] <= 32'h0;
memory[3020] <= 32'h0;
memory[3021] <= 32'h0;
memory[3022] <= 32'h0;
memory[3023] <= 32'h0;
memory[3024] <= 32'h0;
memory[3025] <= 32'h0;
memory[3026] <= 32'h0;
memory[3027] <= 32'h0;
memory[3028] <= 32'h0;
memory[3029] <= 32'h0;
memory[3030] <= 32'h0;
memory[3031] <= 32'h0;
memory[3032] <= 32'h0;
memory[3033] <= 32'h0;
memory[3034] <= 32'h0;
memory[3035] <= 32'h0;
memory[3036] <= 32'h0;
memory[3037] <= 32'h0;
memory[3038] <= 32'h0;
memory[3039] <= 32'h0;
memory[3040] <= 32'h0;
memory[3041] <= 32'h0;
memory[3042] <= 32'h0;
memory[3043] <= 32'h0;
memory[3044] <= 32'h0;
memory[3045] <= 32'h0;
memory[3046] <= 32'h0;
memory[3047] <= 32'h0;
memory[3048] <= 32'h0;
memory[3049] <= 32'h0;
memory[3050] <= 32'h0;
memory[3051] <= 32'h0;
memory[3052] <= 32'h0;
memory[3053] <= 32'h0;
memory[3054] <= 32'h0;
memory[3055] <= 32'h0;
memory[3056] <= 32'h0;
memory[3057] <= 32'h0;
memory[3058] <= 32'h0;
memory[3059] <= 32'h0;
memory[3060] <= 32'h0;
memory[3061] <= 32'h0;
memory[3062] <= 32'h0;
memory[3063] <= 32'h0;
memory[3064] <= 32'h0;
memory[3065] <= 32'h0;
memory[3066] <= 32'h0;
memory[3067] <= 32'h0;
memory[3068] <= 32'h0;
memory[3069] <= 32'h0;
memory[3070] <= 32'h0;
memory[3071] <= 32'h0;
memory[3072] <= 32'h0;
memory[3073] <= 32'h0;
memory[3074] <= 32'h0;
memory[3075] <= 32'h0;
memory[3076] <= 32'h0;
memory[3077] <= 32'h0;
memory[3078] <= 32'h0;
memory[3079] <= 32'h0;
memory[3080] <= 32'h0;
memory[3081] <= 32'h0;
memory[3082] <= 32'h0;
memory[3083] <= 32'h0;
memory[3084] <= 32'h0;
memory[3085] <= 32'h0;
memory[3086] <= 32'h0;
memory[3087] <= 32'h0;
memory[3088] <= 32'h0;
memory[3089] <= 32'h0;
memory[3090] <= 32'h0;
memory[3091] <= 32'h0;
memory[3092] <= 32'h0;
memory[3093] <= 32'h0;
memory[3094] <= 32'h0;
memory[3095] <= 32'h0;
memory[3096] <= 32'h0;
memory[3097] <= 32'h0;
memory[3098] <= 32'h0;
memory[3099] <= 32'h0;
memory[3100] <= 32'h0;
memory[3101] <= 32'h0;
memory[3102] <= 32'h0;
memory[3103] <= 32'h0;
memory[3104] <= 32'h0;
memory[3105] <= 32'h0;
memory[3106] <= 32'h0;
memory[3107] <= 32'h0;
memory[3108] <= 32'h0;
memory[3109] <= 32'h0;
memory[3110] <= 32'h0;
memory[3111] <= 32'h0;
memory[3112] <= 32'h0;
memory[3113] <= 32'h0;
memory[3114] <= 32'h0;
memory[3115] <= 32'h0;
memory[3116] <= 32'h0;
memory[3117] <= 32'h0;
memory[3118] <= 32'h0;
memory[3119] <= 32'h0;
memory[3120] <= 32'h0;
memory[3121] <= 32'h0;
memory[3122] <= 32'h0;
memory[3123] <= 32'h0;
memory[3124] <= 32'h0;
memory[3125] <= 32'h0;
memory[3126] <= 32'h0;
memory[3127] <= 32'h0;
memory[3128] <= 32'h0;
memory[3129] <= 32'h0;
memory[3130] <= 32'h0;
memory[3131] <= 32'h0;
memory[3132] <= 32'h0;
memory[3133] <= 32'h0;
memory[3134] <= 32'h0;
memory[3135] <= 32'h0;
memory[3136] <= 32'h0;
memory[3137] <= 32'h0;
memory[3138] <= 32'h0;
memory[3139] <= 32'h0;
memory[3140] <= 32'h0;
memory[3141] <= 32'h0;
memory[3142] <= 32'h0;
memory[3143] <= 32'h0;
memory[3144] <= 32'h0;
memory[3145] <= 32'h0;
memory[3146] <= 32'h0;
memory[3147] <= 32'h0;
memory[3148] <= 32'h0;
memory[3149] <= 32'h0;
memory[3150] <= 32'h0;
memory[3151] <= 32'h0;
memory[3152] <= 32'h0;
memory[3153] <= 32'h0;
memory[3154] <= 32'h0;
memory[3155] <= 32'h0;
memory[3156] <= 32'h0;
memory[3157] <= 32'h0;
memory[3158] <= 32'h0;
memory[3159] <= 32'h0;
memory[3160] <= 32'h0;
memory[3161] <= 32'h0;
memory[3162] <= 32'h0;
memory[3163] <= 32'h0;
memory[3164] <= 32'h0;
memory[3165] <= 32'h0;
memory[3166] <= 32'h0;
memory[3167] <= 32'h0;
memory[3168] <= 32'h0;
memory[3169] <= 32'h0;
memory[3170] <= 32'h0;
memory[3171] <= 32'h0;
memory[3172] <= 32'h0;
memory[3173] <= 32'h0;
memory[3174] <= 32'h0;
memory[3175] <= 32'h0;
memory[3176] <= 32'h0;
memory[3177] <= 32'h0;
memory[3178] <= 32'h0;
memory[3179] <= 32'h0;
memory[3180] <= 32'h0;
memory[3181] <= 32'h0;
memory[3182] <= 32'h0;
memory[3183] <= 32'h0;
memory[3184] <= 32'h0;
memory[3185] <= 32'h0;
memory[3186] <= 32'h0;
memory[3187] <= 32'h0;
memory[3188] <= 32'h0;
memory[3189] <= 32'h0;
memory[3190] <= 32'h0;
memory[3191] <= 32'h0;
memory[3192] <= 32'h0;
memory[3193] <= 32'h0;
memory[3194] <= 32'h0;
memory[3195] <= 32'h0;
memory[3196] <= 32'h0;
memory[3197] <= 32'h0;
memory[3198] <= 32'h0;
memory[3199] <= 32'h0;
memory[3200] <= 32'h0;
memory[3201] <= 32'h0;
memory[3202] <= 32'h0;
memory[3203] <= 32'h0;
memory[3204] <= 32'h0;
memory[3205] <= 32'h0;
memory[3206] <= 32'h0;
memory[3207] <= 32'h0;
memory[3208] <= 32'h0;
memory[3209] <= 32'h0;
memory[3210] <= 32'h0;
memory[3211] <= 32'h0;
memory[3212] <= 32'h0;
memory[3213] <= 32'h0;
memory[3214] <= 32'h0;
memory[3215] <= 32'h0;
memory[3216] <= 32'h0;
memory[3217] <= 32'h0;
memory[3218] <= 32'h0;
memory[3219] <= 32'h0;
memory[3220] <= 32'h0;
memory[3221] <= 32'h0;
memory[3222] <= 32'h0;
memory[3223] <= 32'h0;
memory[3224] <= 32'h0;
memory[3225] <= 32'h0;
memory[3226] <= 32'h0;
memory[3227] <= 32'h0;
memory[3228] <= 32'h0;
memory[3229] <= 32'h0;
memory[3230] <= 32'h0;
memory[3231] <= 32'h0;
memory[3232] <= 32'h0;
memory[3233] <= 32'h0;
memory[3234] <= 32'h0;
memory[3235] <= 32'h0;
memory[3236] <= 32'h0;
memory[3237] <= 32'h0;
memory[3238] <= 32'h0;
memory[3239] <= 32'h0;
memory[3240] <= 32'h0;
memory[3241] <= 32'h0;
memory[3242] <= 32'h0;
memory[3243] <= 32'h0;
memory[3244] <= 32'h0;
memory[3245] <= 32'h0;
memory[3246] <= 32'h0;
memory[3247] <= 32'h0;
memory[3248] <= 32'h0;
memory[3249] <= 32'h0;
memory[3250] <= 32'h0;
memory[3251] <= 32'h0;
memory[3252] <= 32'h0;
memory[3253] <= 32'h0;
memory[3254] <= 32'h0;
memory[3255] <= 32'h0;
memory[3256] <= 32'h0;
memory[3257] <= 32'h0;
memory[3258] <= 32'h0;
memory[3259] <= 32'h0;
memory[3260] <= 32'h0;
memory[3261] <= 32'h0;
memory[3262] <= 32'h0;
memory[3263] <= 32'h0;
memory[3264] <= 32'h0;
memory[3265] <= 32'h0;
memory[3266] <= 32'h0;
memory[3267] <= 32'h0;
memory[3268] <= 32'h0;
memory[3269] <= 32'h0;
memory[3270] <= 32'h0;
memory[3271] <= 32'h0;
memory[3272] <= 32'h0;
memory[3273] <= 32'h0;
memory[3274] <= 32'h0;
memory[3275] <= 32'h0;
memory[3276] <= 32'h0;
memory[3277] <= 32'h0;
memory[3278] <= 32'h0;
memory[3279] <= 32'h0;
memory[3280] <= 32'h0;
memory[3281] <= 32'h0;
memory[3282] <= 32'h0;
memory[3283] <= 32'h0;
memory[3284] <= 32'h0;
memory[3285] <= 32'h0;
memory[3286] <= 32'h0;
memory[3287] <= 32'h0;
memory[3288] <= 32'h0;
memory[3289] <= 32'h0;
memory[3290] <= 32'h0;
memory[3291] <= 32'h0;
memory[3292] <= 32'h0;
memory[3293] <= 32'h0;
memory[3294] <= 32'h0;
memory[3295] <= 32'h0;
memory[3296] <= 32'h0;
memory[3297] <= 32'h0;
memory[3298] <= 32'h0;
memory[3299] <= 32'h0;
memory[3300] <= 32'h0;
memory[3301] <= 32'h0;
memory[3302] <= 32'h0;
memory[3303] <= 32'h0;
memory[3304] <= 32'h0;
memory[3305] <= 32'h0;
memory[3306] <= 32'h0;
memory[3307] <= 32'h0;
memory[3308] <= 32'h0;
memory[3309] <= 32'h0;
memory[3310] <= 32'h0;
memory[3311] <= 32'h0;
memory[3312] <= 32'h0;
memory[3313] <= 32'h0;
memory[3314] <= 32'h0;
memory[3315] <= 32'h0;
memory[3316] <= 32'h0;
memory[3317] <= 32'h0;
memory[3318] <= 32'h0;
memory[3319] <= 32'h0;
memory[3320] <= 32'h0;
memory[3321] <= 32'h0;
memory[3322] <= 32'h0;
memory[3323] <= 32'h0;
memory[3324] <= 32'h0;
memory[3325] <= 32'h0;
memory[3326] <= 32'h0;
memory[3327] <= 32'h0;
memory[3328] <= 32'h0;
memory[3329] <= 32'h0;
memory[3330] <= 32'h0;
memory[3331] <= 32'h0;
memory[3332] <= 32'h0;
memory[3333] <= 32'h0;
memory[3334] <= 32'h0;
memory[3335] <= 32'h0;
memory[3336] <= 32'h0;
memory[3337] <= 32'h0;
memory[3338] <= 32'h0;
memory[3339] <= 32'h0;
memory[3340] <= 32'h0;
memory[3341] <= 32'h0;
memory[3342] <= 32'h0;
memory[3343] <= 32'h0;
memory[3344] <= 32'h0;
memory[3345] <= 32'h0;
memory[3346] <= 32'h0;
memory[3347] <= 32'h0;
memory[3348] <= 32'h0;
memory[3349] <= 32'h0;
memory[3350] <= 32'h0;
memory[3351] <= 32'h0;
memory[3352] <= 32'h0;
memory[3353] <= 32'h0;
memory[3354] <= 32'h0;
memory[3355] <= 32'h0;
memory[3356] <= 32'h0;
memory[3357] <= 32'h0;
memory[3358] <= 32'h0;
memory[3359] <= 32'h0;
memory[3360] <= 32'h0;
memory[3361] <= 32'h0;
memory[3362] <= 32'h0;
memory[3363] <= 32'h0;
memory[3364] <= 32'h0;
memory[3365] <= 32'h0;
memory[3366] <= 32'h0;
memory[3367] <= 32'h0;
memory[3368] <= 32'h0;
memory[3369] <= 32'h0;
memory[3370] <= 32'h0;
memory[3371] <= 32'h0;
memory[3372] <= 32'h0;
memory[3373] <= 32'h0;
memory[3374] <= 32'h0;
memory[3375] <= 32'h0;
memory[3376] <= 32'h0;
memory[3377] <= 32'h0;
memory[3378] <= 32'h0;
memory[3379] <= 32'h0;
memory[3380] <= 32'h0;
memory[3381] <= 32'h0;
memory[3382] <= 32'h0;
memory[3383] <= 32'h0;
memory[3384] <= 32'h0;
memory[3385] <= 32'h0;
memory[3386] <= 32'h0;
memory[3387] <= 32'h0;
memory[3388] <= 32'h0;
memory[3389] <= 32'h0;
memory[3390] <= 32'h0;
memory[3391] <= 32'h0;
memory[3392] <= 32'h0;
memory[3393] <= 32'h0;
memory[3394] <= 32'h0;
memory[3395] <= 32'h0;
memory[3396] <= 32'h0;
memory[3397] <= 32'h0;
memory[3398] <= 32'h0;
memory[3399] <= 32'h0;
memory[3400] <= 32'h0;
memory[3401] <= 32'h0;
memory[3402] <= 32'h0;
memory[3403] <= 32'h0;
memory[3404] <= 32'h0;
memory[3405] <= 32'h0;
memory[3406] <= 32'h0;
memory[3407] <= 32'h0;
memory[3408] <= 32'h0;
memory[3409] <= 32'h0;
memory[3410] <= 32'h0;
memory[3411] <= 32'h0;
memory[3412] <= 32'h0;
memory[3413] <= 32'h0;
memory[3414] <= 32'h0;
memory[3415] <= 32'h0;
memory[3416] <= 32'h0;
memory[3417] <= 32'h0;
memory[3418] <= 32'h0;
memory[3419] <= 32'h0;
memory[3420] <= 32'h0;
memory[3421] <= 32'h0;
memory[3422] <= 32'h0;
memory[3423] <= 32'h0;
memory[3424] <= 32'h0;
memory[3425] <= 32'h0;
memory[3426] <= 32'h0;
memory[3427] <= 32'h0;
memory[3428] <= 32'h0;
memory[3429] <= 32'h0;
memory[3430] <= 32'h0;
memory[3431] <= 32'h0;
memory[3432] <= 32'h0;
memory[3433] <= 32'h0;
memory[3434] <= 32'h0;
memory[3435] <= 32'h0;
memory[3436] <= 32'h0;
memory[3437] <= 32'h0;
memory[3438] <= 32'h0;
memory[3439] <= 32'h0;
memory[3440] <= 32'h0;
memory[3441] <= 32'h0;
memory[3442] <= 32'h0;
memory[3443] <= 32'h1;
memory[3444] <= 32'h1;
memory[3445] <= 32'h1;
memory[3446] <= 32'h1;
memory[3447] <= 32'h1;
memory[3448] <= 32'h1;
memory[3449] <= 32'h1;
memory[3450] <= 32'h1;
memory[3451] <= 32'h1;
memory[3452] <= 32'h1;
memory[3453] <= 32'h1;
memory[3454] <= 32'h1;
memory[3455] <= 32'h1;
memory[3456] <= 32'h1;
memory[3457] <= 32'h1;
memory[3458] <= 32'h1;
memory[3459] <= 32'h20;
memory[3460] <= 32'h20;
memory[3461] <= 32'h4;
memory[3462] <= 32'h4;
memory[3463] <= 32'h1;
memory[3464] <= 32'h1;
memory[3465] <= 32'h1;
memory[3466] <= 32'h1;
memory[3467] <= 32'h1;
memory[3468] <= 32'h0;
memory[3469] <= 32'h0;
memory[3470] <= 32'h0;
memory[3471] <= 32'h0;
memory[3472] <= 32'h0;
memory[3473] <= 32'h0;
memory[3474] <= 32'h0;
memory[3475] <= 32'h0;
memory[3476] <= 32'h0;
memory[3477] <= 32'h0;
memory[3478] <= 32'h0;
memory[3479] <= 32'h0;
memory[3480] <= 32'h0;
memory[3481] <= 32'h0;
memory[3482] <= 32'h0;
memory[3483] <= 32'h0;
memory[3484] <= 32'h0;
memory[3485] <= 32'h0;
memory[3486] <= 32'h0;
memory[3487] <= 32'h0;
memory[3488] <= 32'h0;
memory[3489] <= 32'h0;
memory[3490] <= 32'h0;
memory[3491] <= 32'h0;
memory[3492] <= 32'h0;
memory[3493] <= 32'h0;
memory[3494] <= 32'h0;
memory[3495] <= 32'h1;
memory[3496] <= 32'h1;
memory[3497] <= 32'h1;
memory[3498] <= 32'h1;
memory[3499] <= 32'h1;
memory[3500] <= 32'h0;
memory[3501] <= 32'h0;
memory[3502] <= 32'h0;
memory[3503] <= 32'h0;
memory[3504] <= 32'h0;
memory[3505] <= 32'h0;
memory[3506] <= 32'h0;
memory[3507] <= 32'h0;
memory[3508] <= 32'h0;
memory[3509] <= 32'h0;
memory[3510] <= 32'h0;
memory[3511] <= 32'h0;
memory[3512] <= 32'h0;
memory[3513] <= 32'h0;
memory[3514] <= 32'h0;
memory[3515] <= 32'h0;
memory[3516] <= 32'h0;
memory[3517] <= 32'h0;
memory[3518] <= 32'h0;
memory[3519] <= 32'h0;
memory[3520] <= 32'h0;
memory[3521] <= 32'h0;
memory[3522] <= 32'h0;
memory[3523] <= 32'h0;
memory[3524] <= 32'h0;
memory[3525] <= 32'h0;
memory[3526] <= 32'h0;
memory[3527] <= 32'h1;
memory[3528] <= 32'h1;
memory[3529] <= 32'h1;
memory[3530] <= 32'h1;
memory[3531] <= 32'h1;
memory[3532] <= 32'h0;
memory[3533] <= 32'h0;
memory[3534] <= 32'h0;
memory[3535] <= 32'h0;
memory[3536] <= 32'h0;
memory[3537] <= 32'h0;
memory[3538] <= 32'h0;
memory[3539] <= 32'h0;
memory[3540] <= 32'h0;
memory[3541] <= 32'h0;
memory[3542] <= 32'h0;
memory[3543] <= 32'h0;
memory[3544] <= 32'h0;
memory[3545] <= 32'h0;
memory[3546] <= 32'h0;
memory[3547] <= 32'h0;
memory[3548] <= 32'h0;
memory[3549] <= 32'h0;
memory[3550] <= 32'h0;
memory[3551] <= 32'h0;
memory[3552] <= 32'h0;
memory[3553] <= 32'h0;
memory[3554] <= 32'h0;
memory[3555] <= 32'h0;
memory[3556] <= 32'h0;
memory[3557] <= 32'h0;
memory[3558] <= 32'h0;
memory[3559] <= 32'h1;
memory[3560] <= 32'h1;
memory[3561] <= 32'h1;
memory[3562] <= 32'h1;
memory[3563] <= 32'h1;
memory[3564] <= 32'h0;
memory[3565] <= 32'h0;
memory[3566] <= 32'h0;
memory[3567] <= 32'h0;
memory[3568] <= 32'h0;
memory[3569] <= 32'h0;
memory[3570] <= 32'h0;
memory[3571] <= 32'h0;
memory[3572] <= 32'h0;
memory[3573] <= 32'h0;
memory[3574] <= 32'h0;
memory[3575] <= 32'h0;
memory[3576] <= 32'h0;
memory[3577] <= 32'h0;
memory[3578] <= 32'h0;
memory[3579] <= 32'h0;
memory[3580] <= 32'h0;
memory[3581] <= 32'h0;
memory[3582] <= 32'h0;
memory[3583] <= 32'h0;
memory[3584] <= 32'h0;
memory[3585] <= 32'h0;
memory[3586] <= 32'h0;
memory[3587] <= 32'h0;
memory[3588] <= 32'h0;
memory[3589] <= 32'h0;
memory[3590] <= 32'h0;
memory[3591] <= 32'h0;
memory[3592] <= 32'h0;
memory[3593] <= 32'h0;
memory[3594] <= 32'h0;
memory[3595] <= 32'h0;
memory[3596] <= 32'h0;
memory[3597] <= 32'h0;
memory[3598] <= 32'h0;
memory[3599] <= 32'h0;
memory[3600] <= 32'h0;
memory[3601] <= 32'h0;
memory[3602] <= 32'h0;
memory[3603] <= 32'h0;
memory[3604] <= 32'h0;
memory[3605] <= 32'h0;
memory[3606] <= 32'h0;
memory[3607] <= 32'h0;
memory[3608] <= 32'h0;
memory[3609] <= 32'h0;
memory[3610] <= 32'h0;
memory[3611] <= 32'h0;
memory[3612] <= 32'h0;
memory[3613] <= 32'h0;
memory[3614] <= 32'h0;
memory[3615] <= 32'h0;
memory[3616] <= 32'h0;
memory[3617] <= 32'h0;
memory[3618] <= 32'h0;
memory[3619] <= 32'h0;
memory[3620] <= 32'h0;
memory[3621] <= 32'h0;
memory[3622] <= 32'h0;
memory[3623] <= 32'h0;
memory[3624] <= 32'h0;
memory[3625] <= 32'h0;
memory[3626] <= 32'h0;
memory[3627] <= 32'h0;
memory[3628] <= 32'h0;
memory[3629] <= 32'h0;
memory[3630] <= 32'h0;
memory[3631] <= 32'h0;
memory[3632] <= 32'h0;
memory[3633] <= 32'h0;
memory[3634] <= 32'h0;
memory[3635] <= 32'h0;
memory[3636] <= 32'h0;
memory[3637] <= 32'h0;
memory[3638] <= 32'h0;
memory[3639] <= 32'h0;
memory[3640] <= 32'h0;
memory[3641] <= 32'h0;
memory[3642] <= 32'h0;
memory[3643] <= 32'h0;
memory[3644] <= 32'h0;
memory[3645] <= 32'h0;
memory[3646] <= 32'h0;
memory[3647] <= 32'h0;
memory[3648] <= 32'h0;
memory[3649] <= 32'h0;
memory[3650] <= 32'h0;
memory[3651] <= 32'h0;
memory[3652] <= 32'h0;
memory[3653] <= 32'h0;
memory[3654] <= 32'h0;
memory[3655] <= 32'h0;
memory[3656] <= 32'h0;
memory[3657] <= 32'h0;
memory[3658] <= 32'h0;
memory[3659] <= 32'h0;
memory[3660] <= 32'h0;
memory[3661] <= 32'h0;
memory[3662] <= 32'h0;
memory[3663] <= 32'h0;
memory[3664] <= 32'h0;
memory[3665] <= 32'h0;
memory[3666] <= 32'h0;
memory[3667] <= 32'h0;
memory[3668] <= 32'h0;
memory[3669] <= 32'h0;
memory[3670] <= 32'h0;
memory[3671] <= 32'h0;
memory[3672] <= 32'h0;
memory[3673] <= 32'h0;
memory[3674] <= 32'h0;
memory[3675] <= 32'h0;
memory[3676] <= 32'h0;
memory[3677] <= 32'h0;
memory[3678] <= 32'h0;
memory[3679] <= 32'h0;
memory[3680] <= 32'h0;
memory[3681] <= 32'h0;
memory[3682] <= 32'h0;
memory[3683] <= 32'h0;
memory[3684] <= 32'h0;
memory[3685] <= 32'h0;
memory[3686] <= 32'h0;
memory[3687] <= 32'h0;
memory[3688] <= 32'h0;
memory[3689] <= 32'h0;
memory[3690] <= 32'h0;
memory[3691] <= 32'h0;
memory[3692] <= 32'h0;
memory[3693] <= 32'h0;
memory[3694] <= 32'h0;
memory[3695] <= 32'h0;
memory[3696] <= 32'h0;
memory[3697] <= 32'h0;
memory[3698] <= 32'h0;
memory[3699] <= 32'h0;
memory[3700] <= 32'h0;
memory[3701] <= 32'h0;
memory[3702] <= 32'h0;
memory[3703] <= 32'h0;
memory[3704] <= 32'h0;
memory[3705] <= 32'h0;
memory[3706] <= 32'h0;
memory[3707] <= 32'h0;
memory[3708] <= 32'h0;
memory[3709] <= 32'h0;
memory[3710] <= 32'h0;
memory[3711] <= 32'h0;
memory[3712] <= 32'h0;
memory[3713] <= 32'h0;
memory[3714] <= 32'h0;
memory[3715] <= 32'h0;
memory[3716] <= 32'h0;
memory[3717] <= 32'h0;
memory[3718] <= 32'h0;
memory[3719] <= 32'h0;
memory[3720] <= 32'h0;
memory[3721] <= 32'h0;
memory[3722] <= 32'h0;
memory[3723] <= 32'h0;
memory[3724] <= 32'h0;
memory[3725] <= 32'h0;
memory[3726] <= 32'h0;
memory[3727] <= 32'h0;
memory[3728] <= 32'h0;
memory[3729] <= 32'h0;
memory[3730] <= 32'h0;
memory[3731] <= 32'h0;
memory[3732] <= 32'h0;
memory[3733] <= 32'h0;
memory[3734] <= 32'h0;
memory[3735] <= 32'h0;
memory[3736] <= 32'h0;
memory[3737] <= 32'h0;
memory[3738] <= 32'h0;
memory[3739] <= 32'h0;
memory[3740] <= 32'h0;
memory[3741] <= 32'h0;
memory[3742] <= 32'h0;
memory[3743] <= 32'h0;
memory[3744] <= 32'h0;
memory[3745] <= 32'h0;
memory[3746] <= 32'h0;
memory[3747] <= 32'h0;
memory[3748] <= 32'h0;
memory[3749] <= 32'h0;
memory[3750] <= 32'h0;
memory[3751] <= 32'h0;
memory[3752] <= 32'h0;
memory[3753] <= 32'h0;
memory[3754] <= 32'h0;
memory[3755] <= 32'h0;
memory[3756] <= 32'h0;
memory[3757] <= 32'h0;
memory[3758] <= 32'h0;
memory[3759] <= 32'h0;
memory[3760] <= 32'h0;
memory[3761] <= 32'h0;
memory[3762] <= 32'h0;
memory[3763] <= 32'h0;
memory[3764] <= 32'h0;
memory[3765] <= 32'h0;
memory[3766] <= 32'h0;
memory[3767] <= 32'h0;
memory[3768] <= 32'h0;
memory[3769] <= 32'h0;
memory[3770] <= 32'h0;
memory[3771] <= 32'h0;
memory[3772] <= 32'h0;
memory[3773] <= 32'h0;
memory[3774] <= 32'h0;
memory[3775] <= 32'h0;
memory[3776] <= 32'h0;
memory[3777] <= 32'h0;
memory[3778] <= 32'h0;
memory[3779] <= 32'h0;
memory[3780] <= 32'h0;
memory[3781] <= 32'h0;
memory[3782] <= 32'h0;
memory[3783] <= 32'h0;
memory[3784] <= 32'h0;
memory[3785] <= 32'h0;
memory[3786] <= 32'h0;
memory[3787] <= 32'h0;
memory[3788] <= 32'h0;
memory[3789] <= 32'h0;
memory[3790] <= 32'h0;
memory[3791] <= 32'h0;
memory[3792] <= 32'h0;
memory[3793] <= 32'h0;
memory[3794] <= 32'h0;
memory[3795] <= 32'h0;
memory[3796] <= 32'h0;
memory[3797] <= 32'h0;
memory[3798] <= 32'h0;
memory[3799] <= 32'h0;
memory[3800] <= 32'h0;
memory[3801] <= 32'h0;
memory[3802] <= 32'h0;
memory[3803] <= 32'h0;
memory[3804] <= 32'h0;
memory[3805] <= 32'h0;
memory[3806] <= 32'h0;
memory[3807] <= 32'h0;
memory[3808] <= 32'h0;
memory[3809] <= 32'h0;
memory[3810] <= 32'h0;
memory[3811] <= 32'h0;
memory[3812] <= 32'h0;
memory[3813] <= 32'h0;
memory[3814] <= 32'h0;
memory[3815] <= 32'h0;
memory[3816] <= 32'h0;
memory[3817] <= 32'h0;
memory[3818] <= 32'h0;
memory[3819] <= 32'h0;
memory[3820] <= 32'h0;
memory[3821] <= 32'h0;
memory[3822] <= 32'h0;
memory[3823] <= 32'h0;
memory[3824] <= 32'h0;
memory[3825] <= 32'h0;
memory[3826] <= 32'h0;
memory[3827] <= 32'h0;
memory[3828] <= 32'h0;
memory[3829] <= 32'h0;
memory[3830] <= 32'h0;
memory[3831] <= 32'h0;
memory[3832] <= 32'h0;
memory[3833] <= 32'h0;
memory[3834] <= 32'h0;
memory[3835] <= 32'h0;
memory[3836] <= 32'h0;
memory[3837] <= 32'h0;
memory[3838] <= 32'h0;
memory[3839] <= 32'h0;
memory[3840] <= 32'h0;
memory[3841] <= 32'h0;
memory[3842] <= 32'h0;
memory[3843] <= 32'h0;
memory[3844] <= 32'h0;
memory[3845] <= 32'h0;
memory[3846] <= 32'h0;
memory[3847] <= 32'h0;
memory[3848] <= 32'h0;
memory[3849] <= 32'h0;
memory[3850] <= 32'h0;
memory[3851] <= 32'h0;
memory[3852] <= 32'h0;
memory[3853] <= 32'h0;
memory[3854] <= 32'h0;
memory[3855] <= 32'h0;
memory[3856] <= 32'h0;
memory[3857] <= 32'h0;
memory[3858] <= 32'h0;
memory[3859] <= 32'h0;
memory[3860] <= 32'h0;
memory[3861] <= 32'h0;
memory[3862] <= 32'h0;
memory[3863] <= 32'h0;
memory[3864] <= 32'h0;
memory[3865] <= 32'h0;
memory[3866] <= 32'h0;
memory[3867] <= 32'h0;
memory[3868] <= 32'h0;
memory[3869] <= 32'h0;
memory[3870] <= 32'h0;
memory[3871] <= 32'h0;
memory[3872] <= 32'h0;
memory[3873] <= 32'h0;
memory[3874] <= 32'h0;
memory[3875] <= 32'h0;
memory[3876] <= 32'h0;
memory[3877] <= 32'h0;
memory[3878] <= 32'h0;
memory[3879] <= 32'h0;
memory[3880] <= 32'h0;
memory[3881] <= 32'h0;
memory[3882] <= 32'h0;
memory[3883] <= 32'h0;
memory[3884] <= 32'h0;
memory[3885] <= 32'h0;
memory[3886] <= 32'h0;
memory[3887] <= 32'h0;
memory[3888] <= 32'h0;
memory[3889] <= 32'h0;
memory[3890] <= 32'h0;
memory[3891] <= 32'h0;
memory[3892] <= 32'h0;
memory[3893] <= 32'h0;
memory[3894] <= 32'h0;
memory[3895] <= 32'h0;
memory[3896] <= 32'h0;
memory[3897] <= 32'h0;
memory[3898] <= 32'h0;
memory[3899] <= 32'h0;
memory[3900] <= 32'h0;
memory[3901] <= 32'h0;
memory[3902] <= 32'h0;
memory[3903] <= 32'h0;
memory[3904] <= 32'h0;
memory[3905] <= 32'h0;
memory[3906] <= 32'h0;
memory[3907] <= 32'h0;
memory[3908] <= 32'h0;
memory[3909] <= 32'h0;
memory[3910] <= 32'h0;
memory[3911] <= 32'h0;
memory[3912] <= 32'h0;
memory[3913] <= 32'h0;
memory[3914] <= 32'h0;
memory[3915] <= 32'h0;
memory[3916] <= 32'h0;
memory[3917] <= 32'h0;
memory[3918] <= 32'h0;
memory[3919] <= 32'h0;
memory[3920] <= 32'h0;
memory[3921] <= 32'h0;
memory[3922] <= 32'h0;
memory[3923] <= 32'h0;
memory[3924] <= 32'h0;
memory[3925] <= 32'h0;
memory[3926] <= 32'h0;
memory[3927] <= 32'h0;
memory[3928] <= 32'h0;
memory[3929] <= 32'h0;
memory[3930] <= 32'h0;
memory[3931] <= 32'h0;
memory[3932] <= 32'h0;
memory[3933] <= 32'h0;
memory[3934] <= 32'h0;
memory[3935] <= 32'h0;
memory[3936] <= 32'h0;
memory[3937] <= 32'h0;
memory[3938] <= 32'h0;
memory[3939] <= 32'h0;
memory[3940] <= 32'h0;
memory[3941] <= 32'h0;
memory[3942] <= 32'h0;
memory[3943] <= 32'h0;
memory[3944] <= 32'h0;
memory[3945] <= 32'h0;
memory[3946] <= 32'h0;
memory[3947] <= 32'h0;
memory[3948] <= 32'h0;
memory[3949] <= 32'h0;
memory[3950] <= 32'h0;
memory[3951] <= 32'h0;
memory[3952] <= 32'h0;
memory[3953] <= 32'h0;
memory[3954] <= 32'h0;
memory[3955] <= 32'h0;
memory[3956] <= 32'h0;
memory[3957] <= 32'h0;
memory[3958] <= 32'h0;
memory[3959] <= 32'h0;
memory[3960] <= 32'h0;
memory[3961] <= 32'h0;
memory[3962] <= 32'h0;
memory[3963] <= 32'h0;
memory[3964] <= 32'h0;
memory[3965] <= 32'h0;
memory[3966] <= 32'h0;
memory[3967] <= 32'h0;
memory[3968] <= 32'h0;
memory[3969] <= 32'h0;
memory[3970] <= 32'h0;
memory[3971] <= 32'h0;
memory[3972] <= 32'h0;
memory[3973] <= 32'h0;
memory[3974] <= 32'h0;
memory[3975] <= 32'h0;
memory[3976] <= 32'h0;
memory[3977] <= 32'h0;
memory[3978] <= 32'h0;
memory[3979] <= 32'h0;
memory[3980] <= 32'h0;
memory[3981] <= 32'h0;
memory[3982] <= 32'h0;
memory[3983] <= 32'h0;
memory[3984] <= 32'h0;
memory[3985] <= 32'h0;
memory[3986] <= 32'h0;
memory[3987] <= 32'h0;
memory[3988] <= 32'h0;
memory[3989] <= 32'h0;
memory[3990] <= 32'h0;
memory[3991] <= 32'h0;
memory[3992] <= 32'h0;
memory[3993] <= 32'h0;
memory[3994] <= 32'h0;
memory[3995] <= 32'h0;
memory[3996] <= 32'h0;
memory[3997] <= 32'h0;
memory[3998] <= 32'h0;
memory[3999] <= 32'h0;
memory[4000] <= 32'h0;
memory[4001] <= 32'h0;
memory[4002] <= 32'h0;
memory[4003] <= 32'h0;
memory[4004] <= 32'h0;
memory[4005] <= 32'h0;
memory[4006] <= 32'h0;
memory[4007] <= 32'h0;
memory[4008] <= 32'h0;
memory[4009] <= 32'h0;
memory[4010] <= 32'h0;
memory[4011] <= 32'h0;
memory[4012] <= 32'h0;
memory[4013] <= 32'h0;
memory[4014] <= 32'h0;
memory[4015] <= 32'h0;
memory[4016] <= 32'h0;
memory[4017] <= 32'h0;
memory[4018] <= 32'h0;
memory[4019] <= 32'h0;
memory[4020] <= 32'h0;
memory[4021] <= 32'h0;
memory[4022] <= 32'h0;
memory[4023] <= 32'h0;
memory[4024] <= 32'h0;
memory[4025] <= 32'h0;
memory[4026] <= 32'h0;
memory[4027] <= 32'h0;
memory[4028] <= 32'h0;
memory[4029] <= 32'h0;
memory[4030] <= 32'h0;
memory[4031] <= 32'h0;
memory[4032] <= 32'h0;
memory[4033] <= 32'h0;
memory[4034] <= 32'h0;
memory[4035] <= 32'h0;
memory[4036] <= 32'h0;
memory[4037] <= 32'h0;
memory[4038] <= 32'h0;
memory[4039] <= 32'h0;
memory[4040] <= 32'h0;
memory[4041] <= 32'h0;
memory[4042] <= 32'h0;
memory[4043] <= 32'h0;
memory[4044] <= 32'h0;
memory[4045] <= 32'h0;
memory[4046] <= 32'h0;
memory[4047] <= 32'h0;
memory[4048] <= 32'h0;
memory[4049] <= 32'h0;
memory[4050] <= 32'h0;
memory[4051] <= 32'h0;
memory[4052] <= 32'h0;
memory[4053] <= 32'h0;
memory[4054] <= 32'h0;
memory[4055] <= 32'h0;
memory[4056] <= 32'h0;
memory[4057] <= 32'h0;
memory[4058] <= 32'h0;
memory[4059] <= 32'h0;
memory[4060] <= 32'h0;
memory[4061] <= 32'h0;
memory[4062] <= 32'h0;
memory[4063] <= 32'h0;
memory[4064] <= 32'h0;
memory[4065] <= 32'h0;
memory[4066] <= 32'h0;
memory[4067] <= 32'h0;
memory[4068] <= 32'h0;
memory[4069] <= 32'h0;
memory[4070] <= 32'h0;
memory[4071] <= 32'h0;
memory[4072] <= 32'h0;
memory[4073] <= 32'h0;
memory[4074] <= 32'h0;
memory[4075] <= 32'h0;
memory[4076] <= 32'h0;
memory[4077] <= 32'h0;
memory[4078] <= 32'h0;
memory[4079] <= 32'h0;
memory[4080] <= 32'h0;
memory[4081] <= 32'h0;
memory[4082] <= 32'h0;
memory[4083] <= 32'h0;
memory[4084] <= 32'h0;
memory[4085] <= 32'h0;
memory[4086] <= 32'h0;
memory[4087] <= 32'h0;
memory[4088] <= 32'h0;
memory[4089] <= 32'h0;
memory[4090] <= 32'h0;
memory[4091] <= 32'h0;
memory[4092] <= 32'h0;
memory[4093] <= 32'h0;
memory[4094] <= 32'h0;
memory[4095] <= 32'h0;
memory[4096] <= 32'h0;
memory[4097] <= 32'h0;
memory[4098] <= 32'h0;
memory[4099] <= 32'h0;
memory[4100] <= 32'h0;
memory[4101] <= 32'h0;
memory[4102] <= 32'h0;
memory[4103] <= 32'h0;
memory[4104] <= 32'h0;
memory[4105] <= 32'h0;
memory[4106] <= 32'h0;
memory[4107] <= 32'h0;
memory[4108] <= 32'h0;
memory[4109] <= 32'h0;
memory[4110] <= 32'h0;
memory[4111] <= 32'h0;
memory[4112] <= 32'h0;
memory[4113] <= 32'h0;
memory[4114] <= 32'h0;
memory[4115] <= 32'h0;
memory[4116] <= 32'h0;
memory[4117] <= 32'h0;
memory[4118] <= 32'h0;
memory[4119] <= 32'h0;
memory[4120] <= 32'h0;
memory[4121] <= 32'h0;
memory[4122] <= 32'h0;
memory[4123] <= 32'h0;
memory[4124] <= 32'h0;
memory[4125] <= 32'h0;
memory[4126] <= 32'h0;
memory[4127] <= 32'h0;
memory[4128] <= 32'h0;
memory[4129] <= 32'h0;
memory[4130] <= 32'h0;
memory[4131] <= 32'h0;
memory[4132] <= 32'h0;
memory[4133] <= 32'h0;
memory[4134] <= 32'h0;
memory[4135] <= 32'h0;
memory[4136] <= 32'h0;
memory[4137] <= 32'h0;
memory[4138] <= 32'h0;
memory[4139] <= 32'h0;
memory[4140] <= 32'h0;
memory[4141] <= 32'h0;
memory[4142] <= 32'h0;
memory[4143] <= 32'h0;
memory[4144] <= 32'h0;
memory[4145] <= 32'h0;
memory[4146] <= 32'h0;
memory[4147] <= 32'h0;
memory[4148] <= 32'h0;
memory[4149] <= 32'h0;
memory[4150] <= 32'h0;
memory[4151] <= 32'h0;
memory[4152] <= 32'h0;
memory[4153] <= 32'h0;
memory[4154] <= 32'h0;
memory[4155] <= 32'h0;
memory[4156] <= 32'h0;
memory[4157] <= 32'h0;
memory[4158] <= 32'h0;
memory[4159] <= 32'h0;
memory[4160] <= 32'h0;
memory[4161] <= 32'h0;
memory[4162] <= 32'h0;
memory[4163] <= 32'h0;
memory[4164] <= 32'h0;
memory[4165] <= 32'h0;
memory[4166] <= 32'h0;
memory[4167] <= 32'h0;
memory[4168] <= 32'h0;
memory[4169] <= 32'h0;
memory[4170] <= 32'h0;
memory[4171] <= 32'h0;
memory[4172] <= 32'h0;
memory[4173] <= 32'h0;
memory[4174] <= 32'h0;
memory[4175] <= 32'h0;
memory[4176] <= 32'h0;
memory[4177] <= 32'h0;
memory[4178] <= 32'h0;
memory[4179] <= 32'h0;
memory[4180] <= 32'h0;
memory[4181] <= 32'h0;
memory[4182] <= 32'h0;
memory[4183] <= 32'h0;
memory[4184] <= 32'h0;
memory[4185] <= 32'h0;
memory[4186] <= 32'h0;
memory[4187] <= 32'h0;
memory[4188] <= 32'h0;
memory[4189] <= 32'h0;
memory[4190] <= 32'h0;
memory[4191] <= 32'h0;
memory[4192] <= 32'h0;
memory[4193] <= 32'h0;
memory[4194] <= 32'h0;
memory[4195] <= 32'h0;
memory[4196] <= 32'h0;
memory[4197] <= 32'h0;
memory[4198] <= 32'h0;
memory[4199] <= 32'h0;
memory[4200] <= 32'h0;
memory[4201] <= 32'h0;
memory[4202] <= 32'h0;
memory[4203] <= 32'h0;
memory[4204] <= 32'h0;
memory[4205] <= 32'h0;
memory[4206] <= 32'h0;
memory[4207] <= 32'h0;
memory[4208] <= 32'h0;
memory[4209] <= 32'h0;
memory[4210] <= 32'h0;
memory[4211] <= 32'h0;
memory[4212] <= 32'h0;
memory[4213] <= 32'h0;
memory[4214] <= 32'h0;
memory[4215] <= 32'h0;
memory[4216] <= 32'h0;
memory[4217] <= 32'h0;
memory[4218] <= 32'h0;
memory[4219] <= 32'h0;
memory[4220] <= 32'h0;
memory[4221] <= 32'h0;
memory[4222] <= 32'h0;
memory[4223] <= 32'h0;
memory[4224] <= 32'h0;
memory[4225] <= 32'h0;
memory[4226] <= 32'h0;
memory[4227] <= 32'h0;
memory[4228] <= 32'h0;
memory[4229] <= 32'h0;
memory[4230] <= 32'h0;
memory[4231] <= 32'h0;
memory[4232] <= 32'h0;
memory[4233] <= 32'h0;
memory[4234] <= 32'h0;
memory[4235] <= 32'h0;
memory[4236] <= 32'h0;
memory[4237] <= 32'h0;
memory[4238] <= 32'h0;
memory[4239] <= 32'h0;
memory[4240] <= 32'h0;
memory[4241] <= 32'h0;
memory[4242] <= 32'h0;
memory[4243] <= 32'h0;
memory[4244] <= 32'h0;
memory[4245] <= 32'h0;
memory[4246] <= 32'h0;
memory[4247] <= 32'h0;
memory[4248] <= 32'h0;
memory[4249] <= 32'h0;
memory[4250] <= 32'h0;
memory[4251] <= 32'h0;
memory[4252] <= 32'h0;
memory[4253] <= 32'h0;
memory[4254] <= 32'h0;
memory[4255] <= 32'h0;
memory[4256] <= 32'h0;
memory[4257] <= 32'h0;
memory[4258] <= 32'h0;
memory[4259] <= 32'h0;
memory[4260] <= 32'h0;
memory[4261] <= 32'h0;
memory[4262] <= 32'h0;
memory[4263] <= 32'h0;
memory[4264] <= 32'h0;
memory[4265] <= 32'h0;
memory[4266] <= 32'h0;
memory[4267] <= 32'h0;
memory[4268] <= 32'h0;
memory[4269] <= 32'h0;
memory[4270] <= 32'h0;
memory[4271] <= 32'h0;
memory[4272] <= 32'h0;
memory[4273] <= 32'h0;
memory[4274] <= 32'h0;
memory[4275] <= 32'h0;
memory[4276] <= 32'h0;
memory[4277] <= 32'h0;
memory[4278] <= 32'h0;
memory[4279] <= 32'h0;
memory[4280] <= 32'h0;
memory[4281] <= 32'h0;
memory[4282] <= 32'h0;
memory[4283] <= 32'h0;
memory[4284] <= 32'h0;
memory[4285] <= 32'h0;
memory[4286] <= 32'h0;
memory[4287] <= 32'h0;
memory[4288] <= 32'h0;
memory[4289] <= 32'h0;
memory[4290] <= 32'h0;
memory[4291] <= 32'h0;
memory[4292] <= 32'h0;
memory[4293] <= 32'h0;
memory[4294] <= 32'h0;
memory[4295] <= 32'h0;
memory[4296] <= 32'h0;
memory[4297] <= 32'h0;
memory[4298] <= 32'h0;
memory[4299] <= 32'h0;
memory[4300] <= 32'h0;
memory[4301] <= 32'h0;
memory[4302] <= 32'h0;
memory[4303] <= 32'h0;
memory[4304] <= 32'h0;
memory[4305] <= 32'h0;
memory[4306] <= 32'h0;
memory[4307] <= 32'h0;
memory[4308] <= 32'h0;
memory[4309] <= 32'h0;
memory[4310] <= 32'h0;
memory[4311] <= 32'h0;
memory[4312] <= 32'h0;
memory[4313] <= 32'h0;
memory[4314] <= 32'h0;
memory[4315] <= 32'h0;
memory[4316] <= 32'h0;
memory[4317] <= 32'h0;
memory[4318] <= 32'h0;
memory[4319] <= 32'h0;
memory[4320] <= 32'h0;
memory[4321] <= 32'h0;
memory[4322] <= 32'h0;
memory[4323] <= 32'h0;
memory[4324] <= 32'h0;
memory[4325] <= 32'h0;
memory[4326] <= 32'h0;
memory[4327] <= 32'h0;
memory[4328] <= 32'h0;
memory[4329] <= 32'h0;
memory[4330] <= 32'h0;
memory[4331] <= 32'h0;
memory[4332] <= 32'h0;
memory[4333] <= 32'h0;
memory[4334] <= 32'h0;
memory[4335] <= 32'h0;
memory[4336] <= 32'h0;
memory[4337] <= 32'h0;
memory[4338] <= 32'h0;
memory[4339] <= 32'h0;
memory[4340] <= 32'h0;
memory[4341] <= 32'h0;
memory[4342] <= 32'h0;
memory[4343] <= 32'h0;
memory[4344] <= 32'h0;
memory[4345] <= 32'h0;
memory[4346] <= 32'h0;
memory[4347] <= 32'h0;
memory[4348] <= 32'h0;
memory[4349] <= 32'h0;
memory[4350] <= 32'h0;
memory[4351] <= 32'h0;
memory[4352] <= 32'h0;
memory[4353] <= 32'h0;
memory[4354] <= 32'h0;
memory[4355] <= 32'h0;
memory[4356] <= 32'h0;
memory[4357] <= 32'h0;
memory[4358] <= 32'h0;
memory[4359] <= 32'h0;
memory[4360] <= 32'h0;
memory[4361] <= 32'h0;
memory[4362] <= 32'h0;
memory[4363] <= 32'h0;
memory[4364] <= 32'h0;
memory[4365] <= 32'h0;
memory[4366] <= 32'h0;
memory[4367] <= 32'h0;
memory[4368] <= 32'h0;
memory[4369] <= 32'h0;
memory[4370] <= 32'h0;
memory[4371] <= 32'h0;
memory[4372] <= 32'h0;
memory[4373] <= 32'h0;
memory[4374] <= 32'h0;
memory[4375] <= 32'h0;
memory[4376] <= 32'h0;
memory[4377] <= 32'h0;
memory[4378] <= 32'h0;
memory[4379] <= 32'h0;
memory[4380] <= 32'h0;
memory[4381] <= 32'h0;
memory[4382] <= 32'h0;
memory[4383] <= 32'h0;
memory[4384] <= 32'h0;
memory[4385] <= 32'h0;
memory[4386] <= 32'h0;
memory[4387] <= 32'h0;
memory[4388] <= 32'h0;
memory[4389] <= 32'h0;
memory[4390] <= 32'h0;
memory[4391] <= 32'h0;
memory[4392] <= 32'h0;
memory[4393] <= 32'h0;
memory[4394] <= 32'h0;
memory[4395] <= 32'h0;
memory[4396] <= 32'h0;
memory[4397] <= 32'h0;
memory[4398] <= 32'h0;
memory[4399] <= 32'h0;
memory[4400] <= 32'h0;
memory[4401] <= 32'h0;
memory[4402] <= 32'h0;
memory[4403] <= 32'h0;
memory[4404] <= 32'h0;
memory[4405] <= 32'h0;
memory[4406] <= 32'h0;
memory[4407] <= 32'h0;
memory[4408] <= 32'h0;
memory[4409] <= 32'h0;
memory[4410] <= 32'h0;
memory[4411] <= 32'h0;
memory[4412] <= 32'h0;
memory[4413] <= 32'h0;
memory[4414] <= 32'h0;
memory[4415] <= 32'h0;
memory[4416] <= 32'h0;
memory[4417] <= 32'h0;
memory[4418] <= 32'h0;
memory[4419] <= 32'h0;
memory[4420] <= 32'h0;
memory[4421] <= 32'h0;
memory[4422] <= 32'h0;
memory[4423] <= 32'h0;
memory[4424] <= 32'h0;
memory[4425] <= 32'h0;
memory[4426] <= 32'h0;
memory[4427] <= 32'h0;
memory[4428] <= 32'h0;
memory[4429] <= 32'h0;
memory[4430] <= 32'h0;
memory[4431] <= 32'h0;
memory[4432] <= 32'h0;
memory[4433] <= 32'h0;
memory[4434] <= 32'h0;
memory[4435] <= 32'h0;
memory[4436] <= 32'h0;
memory[4437] <= 32'h0;
memory[4438] <= 32'h0;
memory[4439] <= 32'h0;
memory[4440] <= 32'h0;
memory[4441] <= 32'h0;
memory[4442] <= 32'h0;
memory[4443] <= 32'h0;
memory[4444] <= 32'h0;
memory[4445] <= 32'h0;
memory[4446] <= 32'h0;
memory[4447] <= 32'h0;
memory[4448] <= 32'h0;
memory[4449] <= 32'h0;
memory[4450] <= 32'h0;
memory[4451] <= 32'h0;
memory[4452] <= 32'h0;
memory[4453] <= 32'h0;
memory[4454] <= 32'h0;
memory[4455] <= 32'h0;
memory[4456] <= 32'h0;
memory[4457] <= 32'h0;
memory[4458] <= 32'h0;
memory[4459] <= 32'h0;
memory[4460] <= 32'h0;
memory[4461] <= 32'h0;
memory[4462] <= 32'h0;
memory[4463] <= 32'h0;
memory[4464] <= 32'h0;
memory[4465] <= 32'h0;
memory[4466] <= 32'h0;
memory[4467] <= 32'h0;
memory[4468] <= 32'h0;
memory[4469] <= 32'h0;
memory[4470] <= 32'h0;
memory[4471] <= 32'h0;
memory[4472] <= 32'h0;
memory[4473] <= 32'h0;
memory[4474] <= 32'h0;
memory[4475] <= 32'h0;
memory[4476] <= 32'h0;
memory[4477] <= 32'h0;
memory[4478] <= 32'h0;
memory[4479] <= 32'h0;
memory[4480] <= 32'h0;
memory[4481] <= 32'h0;
memory[4482] <= 32'h0;
memory[4483] <= 32'h0;
memory[4484] <= 32'h0;
memory[4485] <= 32'h0;
memory[4486] <= 32'h0;
memory[4487] <= 32'h1;
memory[4488] <= 32'h1;
memory[4489] <= 32'h1;
memory[4490] <= 32'h1;
memory[4491] <= 32'h1;
memory[4492] <= 32'h1;
memory[4493] <= 32'h1;
memory[4494] <= 32'h1;
memory[4495] <= 32'h1;
memory[4496] <= 32'h1;
memory[4497] <= 32'h1;
memory[4498] <= 32'h1;
memory[4499] <= 32'h1;
memory[4500] <= 32'h1;
memory[4501] <= 32'h1;
memory[4502] <= 32'h1;
memory[4503] <= 32'h32;
memory[4504] <= 32'h20;
memory[4505] <= 32'h8;
memory[4506] <= 32'h4;
memory[4507] <= 32'h0;
memory[4508] <= 32'h0;
memory[4509] <= 32'h0;
memory[4510] <= 32'h0;
memory[4511] <= 32'h0;
memory[4512] <= 32'h0;
memory[4513] <= 32'h0;
memory[4514] <= 32'h0;
memory[4515] <= 32'h0;
memory[4516] <= 32'h0;
memory[4517] <= 32'h0;
memory[4518] <= 32'h0;
memory[4519] <= 32'h0;
memory[4520] <= 32'h0;
memory[4521] <= 32'h0;
memory[4522] <= 32'h0;
memory[4523] <= 32'h0;
memory[4524] <= 32'h0;
memory[4525] <= 32'h0;
memory[4526] <= 32'h0;
memory[4527] <= 32'h0;
memory[4528] <= 32'h0;
memory[4529] <= 32'h0;
memory[4530] <= 32'h0;
memory[4531] <= 32'h0;
memory[4532] <= 32'h0;
memory[4533] <= 32'h0;
memory[4534] <= 32'h0;
memory[4535] <= 32'h0;
memory[4536] <= 32'h0;
memory[4537] <= 32'h0;
memory[4538] <= 32'h0;
memory[4539] <= 32'h0;
memory[4540] <= 32'h0;
memory[4541] <= 32'h0;
memory[4542] <= 32'h0;
memory[4543] <= 32'h0;
memory[4544] <= 32'h0;
memory[4545] <= 32'h0;
memory[4546] <= 32'h0;
memory[4547] <= 32'h0;
memory[4548] <= 32'h0;
memory[4549] <= 32'h0;
memory[4550] <= 32'h0;
memory[4551] <= 32'h0;
memory[4552] <= 32'h0;
memory[4553] <= 32'h0;
memory[4554] <= 32'h0;
memory[4555] <= 32'h0;
memory[4556] <= 32'h0;
memory[4557] <= 32'h0;
memory[4558] <= 32'h0;
memory[4559] <= 32'h0;
memory[4560] <= 32'h0;
memory[4561] <= 32'h0;
memory[4562] <= 32'h0;
memory[4563] <= 32'h0;
memory[4564] <= 32'h0;
memory[4565] <= 32'h0;
memory[4566] <= 32'h0;
memory[4567] <= 32'h0;
memory[4568] <= 32'h0;
memory[4569] <= 32'h0;
memory[4570] <= 32'h0;
memory[4571] <= 32'h0;
memory[4572] <= 32'h0;
memory[4573] <= 32'h0;
memory[4574] <= 32'h0;
memory[4575] <= 32'h0;
memory[4576] <= 32'h0;
memory[4577] <= 32'h0;
memory[4578] <= 32'h0;
memory[4579] <= 32'h0;
memory[4580] <= 32'h0;
memory[4581] <= 32'h0;
memory[4582] <= 32'h0;
memory[4583] <= 32'h0;
memory[4584] <= 32'h0;
memory[4585] <= 32'h0;
memory[4586] <= 32'h0;
memory[4587] <= 32'h0;
memory[4588] <= 32'h0;
memory[4589] <= 32'h0;
memory[4590] <= 32'h0;
memory[4591] <= 32'h0;
memory[4592] <= 32'h0;
memory[4593] <= 32'h0;
memory[4594] <= 32'h0;
memory[4595] <= 32'h0;
memory[4596] <= 32'h0;
memory[4597] <= 32'h0;
memory[4598] <= 32'h0;
memory[4599] <= 32'h0;
memory[4600] <= 32'h0;
memory[4601] <= 32'h0;
memory[4602] <= 32'h0;
memory[4603] <= 32'h0;
memory[4604] <= 32'h0;
memory[4605] <= 32'h0;
memory[4606] <= 32'h0;
memory[4607] <= 32'h0;
memory[4608] <= 32'h0;
memory[4609] <= 32'h0;
memory[4610] <= 32'h0;
memory[4611] <= 32'h0;
memory[4612] <= 32'h0;
memory[4613] <= 32'h0;
memory[4614] <= 32'h0;
memory[4615] <= 32'h0;
memory[4616] <= 32'h0;
memory[4617] <= 32'h0;
memory[4618] <= 32'h0;
memory[4619] <= 32'h0;
memory[4620] <= 32'h0;
memory[4621] <= 32'h0;
memory[4622] <= 32'h0;
memory[4623] <= 32'h0;
memory[4624] <= 32'h0;
memory[4625] <= 32'h0;
memory[4626] <= 32'h0;
memory[4627] <= 32'h0;
memory[4628] <= 32'h0;
memory[4629] <= 32'h0;
memory[4630] <= 32'h0;
memory[4631] <= 32'h0;
memory[4632] <= 32'h0;
memory[4633] <= 32'h0;
memory[4634] <= 32'h0;
memory[4635] <= 32'h0;
memory[4636] <= 32'h0;
memory[4637] <= 32'h0;
memory[4638] <= 32'h0;
memory[4639] <= 32'h0;
memory[4640] <= 32'h0;
memory[4641] <= 32'h0;
memory[4642] <= 32'h0;
memory[4643] <= 32'h0;
memory[4644] <= 32'h0;
memory[4645] <= 32'h0;
memory[4646] <= 32'h0;
memory[4647] <= 32'h0;
memory[4648] <= 32'h0;
memory[4649] <= 32'h0;
memory[4650] <= 32'h0;
memory[4651] <= 32'h0;
memory[4652] <= 32'h0;
memory[4653] <= 32'h0;
memory[4654] <= 32'h0;
memory[4655] <= 32'h0;
memory[4656] <= 32'h0;
memory[4657] <= 32'h0;
memory[4658] <= 32'h0;
memory[4659] <= 32'h0;
memory[4660] <= 32'h0;
memory[4661] <= 32'h0;
memory[4662] <= 32'h0;
memory[4663] <= 32'h0;
memory[4664] <= 32'h0;
memory[4665] <= 32'h0;
memory[4666] <= 32'h0;
memory[4667] <= 32'h0;
memory[4668] <= 32'h0;
memory[4669] <= 32'h0;
memory[4670] <= 32'h0;
memory[4671] <= 32'h0;
memory[4672] <= 32'h0;
memory[4673] <= 32'h0;
memory[4674] <= 32'h0;
memory[4675] <= 32'h0;
memory[4676] <= 32'h0;
memory[4677] <= 32'h0;
memory[4678] <= 32'h0;
memory[4679] <= 32'h0;
memory[4680] <= 32'h0;
memory[4681] <= 32'h0;
memory[4682] <= 32'h0;
memory[4683] <= 32'h0;
memory[4684] <= 32'h0;
memory[4685] <= 32'h0;
memory[4686] <= 32'h0;
memory[4687] <= 32'h0;
memory[4688] <= 32'h0;
memory[4689] <= 32'h0;
memory[4690] <= 32'h0;
memory[4691] <= 32'h0;
memory[4692] <= 32'h0;
memory[4693] <= 32'h0;
memory[4694] <= 32'h0;
memory[4695] <= 32'h0;
memory[4696] <= 32'h0;
memory[4697] <= 32'h0;
memory[4698] <= 32'h0;
memory[4699] <= 32'h0;
memory[4700] <= 32'h0;
memory[4701] <= 32'h0;
memory[4702] <= 32'h0;
memory[4703] <= 32'h0;
memory[4704] <= 32'h0;
memory[4705] <= 32'h0;
memory[4706] <= 32'h0;
memory[4707] <= 32'h0;
memory[4708] <= 32'h0;
memory[4709] <= 32'h0;
memory[4710] <= 32'h0;
memory[4711] <= 32'h0;
memory[4712] <= 32'h0;
memory[4713] <= 32'h0;
memory[4714] <= 32'h0;
memory[4715] <= 32'h0;
memory[4716] <= 32'h0;
memory[4717] <= 32'h0;
memory[4718] <= 32'h0;
memory[4719] <= 32'h0;
memory[4720] <= 32'h0;
memory[4721] <= 32'h0;
memory[4722] <= 32'h0;
memory[4723] <= 32'h0;
memory[4724] <= 32'h0;
memory[4725] <= 32'h0;
memory[4726] <= 32'h0;
memory[4727] <= 32'h0;
memory[4728] <= 32'h0;
memory[4729] <= 32'h0;
memory[4730] <= 32'h0;
memory[4731] <= 32'h0;
memory[4732] <= 32'h0;
memory[4733] <= 32'h0;
memory[4734] <= 32'h0;
memory[4735] <= 32'h0;
memory[4736] <= 32'h0;
memory[4737] <= 32'h0;
memory[4738] <= 32'h0;
memory[4739] <= 32'h0;
memory[4740] <= 32'h0;
memory[4741] <= 32'h0;
memory[4742] <= 32'h0;
memory[4743] <= 32'h0;
memory[4744] <= 32'h0;
memory[4745] <= 32'h0;
memory[4746] <= 32'h0;
memory[4747] <= 32'h0;
memory[4748] <= 32'h0;
memory[4749] <= 32'h0;
memory[4750] <= 32'h0;
memory[4751] <= 32'h0;
memory[4752] <= 32'h0;
memory[4753] <= 32'h0;
memory[4754] <= 32'h0;
memory[4755] <= 32'h0;
memory[4756] <= 32'h0;
memory[4757] <= 32'h0;
memory[4758] <= 32'h0;
memory[4759] <= 32'h0;
memory[4760] <= 32'h0;
memory[4761] <= 32'h0;
memory[4762] <= 32'h0;
memory[4763] <= 32'h0;
memory[4764] <= 32'h0;
memory[4765] <= 32'h0;
memory[4766] <= 32'h0;
memory[4767] <= 32'h0;
memory[4768] <= 32'h0;
memory[4769] <= 32'h0;
memory[4770] <= 32'h0;
memory[4771] <= 32'h0;
memory[4772] <= 32'h0;
memory[4773] <= 32'h0;
memory[4774] <= 32'h0;
memory[4775] <= 32'h0;
memory[4776] <= 32'h0;
memory[4777] <= 32'h0;
memory[4778] <= 32'h0;
memory[4779] <= 32'h0;
memory[4780] <= 32'h0;
memory[4781] <= 32'h0;
memory[4782] <= 32'h0;
memory[4783] <= 32'h0;
memory[4784] <= 32'h0;
memory[4785] <= 32'h0;
memory[4786] <= 32'h0;
memory[4787] <= 32'h0;
memory[4788] <= 32'h0;
memory[4789] <= 32'h0;
memory[4790] <= 32'h0;
memory[4791] <= 32'h0;
memory[4792] <= 32'h0;
memory[4793] <= 32'h0;
memory[4794] <= 32'h0;
memory[4795] <= 32'h0;
memory[4796] <= 32'h0;
memory[4797] <= 32'h0;
memory[4798] <= 32'h0;
memory[4799] <= 32'h0;
memory[4800] <= 32'h0;
memory[4801] <= 32'h0;
memory[4802] <= 32'h0;
memory[4803] <= 32'h0;
memory[4804] <= 32'h0;
memory[4805] <= 32'h0;
memory[4806] <= 32'h0;
memory[4807] <= 32'h0;
memory[4808] <= 32'h0;
memory[4809] <= 32'h0;
memory[4810] <= 32'h0;
memory[4811] <= 32'h0;
memory[4812] <= 32'h0;
memory[4813] <= 32'h0;
memory[4814] <= 32'h0;
memory[4815] <= 32'h0;
memory[4816] <= 32'h0;
memory[4817] <= 32'h0;
memory[4818] <= 32'h0;
memory[4819] <= 32'h0;
memory[4820] <= 32'h0;
memory[4821] <= 32'h0;
memory[4822] <= 32'h0;
memory[4823] <= 32'h0;
memory[4824] <= 32'h0;
memory[4825] <= 32'h0;
memory[4826] <= 32'h0;
memory[4827] <= 32'h0;
memory[4828] <= 32'h0;
memory[4829] <= 32'h0;
memory[4830] <= 32'h0;
memory[4831] <= 32'h0;
memory[4832] <= 32'h0;
memory[4833] <= 32'h0;
memory[4834] <= 32'h0;
memory[4835] <= 32'h0;
memory[4836] <= 32'h0;
memory[4837] <= 32'h0;
memory[4838] <= 32'h0;
memory[4839] <= 32'h0;
memory[4840] <= 32'h0;
memory[4841] <= 32'h0;
memory[4842] <= 32'h0;
memory[4843] <= 32'h0;
memory[4844] <= 32'h0;
memory[4845] <= 32'h0;
memory[4846] <= 32'h0;
memory[4847] <= 32'h0;
memory[4848] <= 32'h0;
memory[4849] <= 32'h0;
memory[4850] <= 32'h0;
memory[4851] <= 32'h0;
memory[4852] <= 32'h0;
memory[4853] <= 32'h0;
memory[4854] <= 32'h0;
memory[4855] <= 32'h0;
memory[4856] <= 32'h0;
memory[4857] <= 32'h0;
memory[4858] <= 32'h0;
memory[4859] <= 32'h0;
memory[4860] <= 32'h0;
memory[4861] <= 32'h0;
memory[4862] <= 32'h0;
memory[4863] <= 32'h0;
memory[4864] <= 32'h0;
memory[4865] <= 32'h0;
memory[4866] <= 32'h0;
memory[4867] <= 32'h0;
memory[4868] <= 32'h0;
memory[4869] <= 32'h0;
memory[4870] <= 32'h0;
memory[4871] <= 32'h0;
memory[4872] <= 32'h0;
memory[4873] <= 32'h0;
memory[4874] <= 32'h0;
memory[4875] <= 32'h0;
memory[4876] <= 32'h0;
memory[4877] <= 32'h0;
memory[4878] <= 32'h0;
memory[4879] <= 32'h0;
memory[4880] <= 32'h0;
memory[4881] <= 32'h0;
memory[4882] <= 32'h0;
memory[4883] <= 32'h0;
memory[4884] <= 32'h0;
memory[4885] <= 32'h0;
memory[4886] <= 32'h0;
memory[4887] <= 32'h0;
memory[4888] <= 32'h0;
memory[4889] <= 32'h0;
memory[4890] <= 32'h0;
memory[4891] <= 32'h0;
memory[4892] <= 32'h0;
memory[4893] <= 32'h0;
memory[4894] <= 32'h0;
memory[4895] <= 32'h0;
memory[4896] <= 32'h0;
memory[4897] <= 32'h0;
memory[4898] <= 32'h0;
memory[4899] <= 32'h0;
memory[4900] <= 32'h0;
memory[4901] <= 32'h0;
memory[4902] <= 32'h0;
memory[4903] <= 32'h0;
memory[4904] <= 32'h0;
memory[4905] <= 32'h0;
memory[4906] <= 32'h0;
memory[4907] <= 32'h0;
memory[4908] <= 32'h0;
memory[4909] <= 32'h0;
memory[4910] <= 32'h0;
memory[4911] <= 32'h0;
memory[4912] <= 32'h0;
memory[4913] <= 32'h0;
memory[4914] <= 32'h0;
memory[4915] <= 32'h0;
memory[4916] <= 32'h0;
memory[4917] <= 32'h0;
memory[4918] <= 32'h0;
memory[4919] <= 32'h0;
memory[4920] <= 32'h0;
memory[4921] <= 32'h0;
memory[4922] <= 32'h0;
memory[4923] <= 32'h0;
memory[4924] <= 32'h0;
memory[4925] <= 32'h0;
memory[4926] <= 32'h0;
memory[4927] <= 32'h0;
memory[4928] <= 32'h0;
memory[4929] <= 32'h0;
memory[4930] <= 32'h0;
memory[4931] <= 32'h0;
memory[4932] <= 32'h0;
memory[4933] <= 32'h0;
memory[4934] <= 32'h0;
memory[4935] <= 32'h0;
memory[4936] <= 32'h0;
memory[4937] <= 32'h0;
memory[4938] <= 32'h0;
memory[4939] <= 32'h0;
memory[4940] <= 32'h0;
memory[4941] <= 32'h0;
memory[4942] <= 32'h0;
memory[4943] <= 32'h0;
memory[4944] <= 32'h0;
memory[4945] <= 32'h0;
memory[4946] <= 32'h0;
memory[4947] <= 32'h0;
memory[4948] <= 32'h0;
memory[4949] <= 32'h0;
memory[4950] <= 32'h0;
memory[4951] <= 32'h0;
memory[4952] <= 32'h0;
memory[4953] <= 32'h0;
memory[4954] <= 32'h0;
memory[4955] <= 32'h0;
memory[4956] <= 32'h0;
memory[4957] <= 32'h0;
memory[4958] <= 32'h0;
memory[4959] <= 32'h0;
memory[4960] <= 32'h0;
memory[4961] <= 32'h0;
memory[4962] <= 32'h0;
memory[4963] <= 32'h0;
memory[4964] <= 32'h0;
memory[4965] <= 32'h0;
memory[4966] <= 32'h0;
memory[4967] <= 32'h0;
memory[4968] <= 32'h0;
memory[4969] <= 32'h0;
memory[4970] <= 32'h0;
memory[4971] <= 32'h0;
memory[4972] <= 32'h0;
memory[4973] <= 32'h0;
memory[4974] <= 32'h0;
memory[4975] <= 32'h0;
memory[4976] <= 32'h0;
memory[4977] <= 32'h0;
memory[4978] <= 32'h0;
memory[4979] <= 32'h0;
memory[4980] <= 32'h0;
memory[4981] <= 32'h0;
memory[4982] <= 32'h0;
memory[4983] <= 32'h0;
memory[4984] <= 32'h0;
memory[4985] <= 32'h0;
memory[4986] <= 32'h0;
memory[4987] <= 32'h0;
memory[4988] <= 32'h0;
memory[4989] <= 32'h0;
memory[4990] <= 32'h0;
memory[4991] <= 32'h0;
memory[4992] <= 32'h0;
memory[4993] <= 32'h0;
memory[4994] <= 32'h0;
memory[4995] <= 32'h0;
memory[4996] <= 32'h0;
memory[4997] <= 32'h0;
memory[4998] <= 32'h0;
memory[4999] <= 32'h0;
memory[5000] <= 32'h0;
memory[5001] <= 32'h0;
memory[5002] <= 32'h0;
memory[5003] <= 32'h0;
memory[5004] <= 32'h0;
memory[5005] <= 32'h0;
memory[5006] <= 32'h0;
memory[5007] <= 32'h0;
memory[5008] <= 32'h0;
memory[5009] <= 32'h0;
memory[5010] <= 32'h0;
memory[5011] <= 32'h0;
memory[5012] <= 32'h0;
memory[5013] <= 32'h0;
memory[5014] <= 32'h0;
memory[5015] <= 32'h0;
memory[5016] <= 32'h0;
memory[5017] <= 32'h0;
memory[5018] <= 32'h0;
memory[5019] <= 32'h0;
memory[5020] <= 32'h0;
memory[5021] <= 32'h0;
memory[5022] <= 32'h0;
memory[5023] <= 32'h0;
memory[5024] <= 32'h0;
memory[5025] <= 32'h0;
memory[5026] <= 32'h0;
memory[5027] <= 32'h0;
memory[5028] <= 32'h0;
memory[5029] <= 32'h0;
memory[5030] <= 32'h0;
memory[5031] <= 32'h0;
memory[5032] <= 32'h0;
memory[5033] <= 32'h0;
memory[5034] <= 32'h0;
memory[5035] <= 32'h0;
memory[5036] <= 32'h0;
memory[5037] <= 32'h0;
memory[5038] <= 32'h0;
memory[5039] <= 32'h0;
memory[5040] <= 32'h0;
memory[5041] <= 32'h0;
memory[5042] <= 32'h0;
memory[5043] <= 32'h0;
memory[5044] <= 32'h0;
memory[5045] <= 32'h0;
memory[5046] <= 32'h0;
memory[5047] <= 32'h0;
memory[5048] <= 32'h0;
memory[5049] <= 32'h0;
memory[5050] <= 32'h0;
memory[5051] <= 32'h0;
memory[5052] <= 32'h0;
memory[5053] <= 32'h0;
memory[5054] <= 32'h0;
memory[5055] <= 32'h0;
memory[5056] <= 32'h0;
memory[5057] <= 32'h0;
memory[5058] <= 32'h0;
memory[5059] <= 32'h0;
memory[5060] <= 32'h0;
memory[5061] <= 32'h0;
memory[5062] <= 32'h0;
memory[5063] <= 32'h0;
memory[5064] <= 32'h0;
memory[5065] <= 32'h0;
memory[5066] <= 32'h0;
memory[5067] <= 32'h0;
memory[5068] <= 32'h0;
memory[5069] <= 32'h0;
memory[5070] <= 32'h0;
memory[5071] <= 32'h0;
memory[5072] <= 32'h0;
memory[5073] <= 32'h0;
memory[5074] <= 32'h0;
memory[5075] <= 32'h0;
memory[5076] <= 32'h0;
memory[5077] <= 32'h0;
memory[5078] <= 32'h0;
memory[5079] <= 32'h0;
memory[5080] <= 32'h0;
memory[5081] <= 32'h0;
memory[5082] <= 32'h0;
memory[5083] <= 32'h0;
memory[5084] <= 32'h0;
memory[5085] <= 32'h0;
memory[5086] <= 32'h0;
memory[5087] <= 32'h0;
memory[5088] <= 32'h0;
memory[5089] <= 32'h0;
memory[5090] <= 32'h0;
memory[5091] <= 32'h0;
memory[5092] <= 32'h0;
memory[5093] <= 32'h0;
memory[5094] <= 32'h0;
memory[5095] <= 32'h0;
memory[5096] <= 32'h0;
memory[5097] <= 32'h0;
memory[5098] <= 32'h0;
memory[5099] <= 32'h0;
memory[5100] <= 32'h0;
memory[5101] <= 32'h0;
memory[5102] <= 32'h0;
memory[5103] <= 32'h0;
memory[5104] <= 32'h0;
memory[5105] <= 32'h0;
memory[5106] <= 32'h0;
memory[5107] <= 32'h0;
memory[5108] <= 32'h0;
memory[5109] <= 32'h0;
memory[5110] <= 32'h0;
memory[5111] <= 32'h0;
memory[5112] <= 32'h0;
memory[5113] <= 32'h0;
memory[5114] <= 32'h0;
memory[5115] <= 32'h0;
memory[5116] <= 32'h0;
memory[5117] <= 32'h0;
memory[5118] <= 32'h0;
memory[5119] <= 32'h0;
memory[5120] <= 32'h0;
memory[5121] <= 32'h0;
memory[5122] <= 32'h0;
memory[5123] <= 32'h0;
memory[5124] <= 32'h0;
memory[5125] <= 32'h0;
memory[5126] <= 32'h0;
memory[5127] <= 32'h0;
memory[5128] <= 32'h0;
memory[5129] <= 32'h0;
memory[5130] <= 32'h0;
memory[5131] <= 32'h0;
memory[5132] <= 32'h0;
memory[5133] <= 32'h0;
memory[5134] <= 32'h0;
memory[5135] <= 32'h0;
memory[5136] <= 32'h0;
memory[5137] <= 32'h0;
memory[5138] <= 32'h0;
memory[5139] <= 32'h0;
memory[5140] <= 32'h0;
memory[5141] <= 32'h0;
memory[5142] <= 32'h0;
memory[5143] <= 32'h0;
memory[5144] <= 32'h0;
memory[5145] <= 32'h0;
memory[5146] <= 32'h0;
memory[5147] <= 32'h0;
memory[5148] <= 32'h0;
memory[5149] <= 32'h0;
memory[5150] <= 32'h0;
memory[5151] <= 32'h0;
memory[5152] <= 32'h0;
memory[5153] <= 32'h0;
memory[5154] <= 32'h0;
memory[5155] <= 32'h0;
memory[5156] <= 32'h0;
memory[5157] <= 32'h0;
memory[5158] <= 32'h0;
memory[5159] <= 32'h0;
memory[5160] <= 32'h0;
memory[5161] <= 32'h0;
memory[5162] <= 32'h0;
memory[5163] <= 32'h0;
memory[5164] <= 32'h0;
memory[5165] <= 32'h0;
memory[5166] <= 32'h0;
memory[5167] <= 32'h0;
memory[5168] <= 32'h0;
memory[5169] <= 32'h0;
memory[5170] <= 32'h0;
memory[5171] <= 32'h0;
memory[5172] <= 32'h0;
memory[5173] <= 32'h0;
memory[5174] <= 32'h0;
memory[5175] <= 32'h0;
memory[5176] <= 32'h0;
memory[5177] <= 32'h0;
memory[5178] <= 32'h0;
memory[5179] <= 32'h0;
memory[5180] <= 32'h0;
memory[5181] <= 32'h0;
memory[5182] <= 32'h0;
memory[5183] <= 32'h0;
memory[5184] <= 32'h0;
memory[5185] <= 32'h0;
memory[5186] <= 32'h0;
memory[5187] <= 32'h0;
memory[5188] <= 32'h0;
memory[5189] <= 32'h0;
memory[5190] <= 32'h0;
memory[5191] <= 32'h0;
memory[5192] <= 32'h0;
memory[5193] <= 32'h0;
memory[5194] <= 32'h0;
memory[5195] <= 32'h0;
memory[5196] <= 32'h0;
memory[5197] <= 32'h0;
memory[5198] <= 32'h0;
memory[5199] <= 32'h0;
memory[5200] <= 32'h0;
memory[5201] <= 32'h0;
memory[5202] <= 32'h0;
memory[5203] <= 32'h0;
memory[5204] <= 32'h0;
memory[5205] <= 32'h0;
memory[5206] <= 32'h0;
memory[5207] <= 32'h0;
memory[5208] <= 32'h0;
memory[5209] <= 32'h0;
memory[5210] <= 32'h0;
memory[5211] <= 32'h0;
memory[5212] <= 32'h0;
memory[5213] <= 32'h0;
memory[5214] <= 32'h0;
memory[5215] <= 32'h0;
memory[5216] <= 32'h0;
memory[5217] <= 32'h0;
memory[5218] <= 32'h0;
memory[5219] <= 32'h0;
memory[5220] <= 32'h0;
memory[5221] <= 32'h0;
memory[5222] <= 32'h0;
memory[5223] <= 32'h0;
memory[5224] <= 32'h0;
memory[5225] <= 32'h0;
memory[5226] <= 32'h0;
memory[5227] <= 32'h0;
memory[5228] <= 32'h0;
memory[5229] <= 32'h0;
memory[5230] <= 32'h0;
memory[5231] <= 32'h0;
memory[5232] <= 32'h0;
memory[5233] <= 32'h0;
memory[5234] <= 32'h0;
memory[5235] <= 32'h0;
memory[5236] <= 32'h0;
memory[5237] <= 32'h0;
memory[5238] <= 32'h0;
memory[5239] <= 32'h0;
memory[5240] <= 32'h0;
memory[5241] <= 32'h0;
memory[5242] <= 32'h0;
memory[5243] <= 32'h0;
memory[5244] <= 32'h0;
memory[5245] <= 32'h0;
memory[5246] <= 32'h0;
memory[5247] <= 32'h0;
memory[5248] <= 32'h0;
memory[5249] <= 32'h0;
memory[5250] <= 32'h0;
memory[5251] <= 32'h0;
memory[5252] <= 32'h0;
memory[5253] <= 32'h0;
memory[5254] <= 32'h0;
memory[5255] <= 32'h0;
memory[5256] <= 32'h0;
memory[5257] <= 32'h0;
memory[5258] <= 32'h0;
memory[5259] <= 32'h0;
memory[5260] <= 32'h0;
memory[5261] <= 32'h0;
memory[5262] <= 32'h0;
memory[5263] <= 32'h0;
memory[5264] <= 32'h0;
memory[5265] <= 32'h0;
memory[5266] <= 32'h0;
memory[5267] <= 32'h0;
memory[5268] <= 32'h0;
memory[5269] <= 32'h0;
memory[5270] <= 32'h0;
memory[5271] <= 32'h0;
memory[5272] <= 32'h0;
memory[5273] <= 32'h0;
memory[5274] <= 32'h0;
memory[5275] <= 32'h0;
memory[5276] <= 32'h0;
memory[5277] <= 32'h0;
memory[5278] <= 32'h0;
memory[5279] <= 32'h0;
memory[5280] <= 32'h0;
memory[5281] <= 32'h0;
memory[5282] <= 32'h0;
memory[5283] <= 32'h0;
memory[5284] <= 32'h0;
memory[5285] <= 32'h0;
memory[5286] <= 32'h0;
memory[5287] <= 32'h0;
memory[5288] <= 32'h0;
memory[5289] <= 32'h0;
memory[5290] <= 32'h0;
memory[5291] <= 32'h0;
memory[5292] <= 32'h0;
memory[5293] <= 32'h0;
memory[5294] <= 32'h0;
memory[5295] <= 32'h0;
memory[5296] <= 32'h0;
memory[5297] <= 32'h0;
memory[5298] <= 32'h0;
memory[5299] <= 32'h0;
memory[5300] <= 32'h0;
memory[5301] <= 32'h0;
memory[5302] <= 32'h0;
memory[5303] <= 32'h0;
memory[5304] <= 32'h0;
memory[5305] <= 32'h0;
memory[5306] <= 32'h0;
memory[5307] <= 32'h0;
memory[5308] <= 32'h0;
memory[5309] <= 32'h0;
memory[5310] <= 32'h0;
memory[5311] <= 32'h0;
memory[5312] <= 32'h0;
memory[5313] <= 32'h0;
memory[5314] <= 32'h0;
memory[5315] <= 32'h0;
memory[5316] <= 32'h0;
memory[5317] <= 32'h0;
memory[5318] <= 32'h0;
memory[5319] <= 32'h0;
memory[5320] <= 32'h0;
memory[5321] <= 32'h0;
memory[5322] <= 32'h0;
memory[5323] <= 32'h0;
memory[5324] <= 32'h0;
memory[5325] <= 32'h0;
memory[5326] <= 32'h0;
memory[5327] <= 32'h0;
memory[5328] <= 32'h0;
memory[5329] <= 32'h0;
memory[5330] <= 32'h0;
memory[5331] <= 32'h0;
memory[5332] <= 32'h0;
memory[5333] <= 32'h0;
memory[5334] <= 32'h0;
memory[5335] <= 32'h0;
memory[5336] <= 32'h0;
memory[5337] <= 32'h0;
memory[5338] <= 32'h0;
memory[5339] <= 32'h0;
memory[5340] <= 32'h0;
memory[5341] <= 32'h0;
memory[5342] <= 32'h0;
memory[5343] <= 32'h0;
memory[5344] <= 32'h0;
memory[5345] <= 32'h0;
memory[5346] <= 32'h0;
memory[5347] <= 32'h0;
memory[5348] <= 32'h0;
memory[5349] <= 32'h0;
memory[5350] <= 32'h0;
memory[5351] <= 32'h0;
memory[5352] <= 32'h0;
memory[5353] <= 32'h0;
memory[5354] <= 32'h0;
memory[5355] <= 32'h0;
memory[5356] <= 32'h0;
memory[5357] <= 32'h0;
memory[5358] <= 32'h0;
memory[5359] <= 32'h0;
memory[5360] <= 32'h0;
memory[5361] <= 32'h0;
memory[5362] <= 32'h0;
memory[5363] <= 32'h0;
memory[5364] <= 32'h0;
memory[5365] <= 32'h0;
memory[5366] <= 32'h0;
memory[5367] <= 32'h0;
memory[5368] <= 32'h0;
memory[5369] <= 32'h0;
memory[5370] <= 32'h0;
memory[5371] <= 32'h0;
memory[5372] <= 32'h0;
memory[5373] <= 32'h0;
memory[5374] <= 32'h0;
memory[5375] <= 32'h0;
memory[5376] <= 32'h0;
memory[5377] <= 32'h0;
memory[5378] <= 32'h0;
memory[5379] <= 32'h0;
memory[5380] <= 32'h0;
memory[5381] <= 32'h0;
memory[5382] <= 32'h0;
memory[5383] <= 32'h0;
memory[5384] <= 32'h0;
memory[5385] <= 32'h0;
memory[5386] <= 32'h0;
memory[5387] <= 32'h0;
memory[5388] <= 32'h0;
memory[5389] <= 32'h0;
memory[5390] <= 32'h0;
memory[5391] <= 32'h0;
memory[5392] <= 32'h0;
memory[5393] <= 32'h0;
memory[5394] <= 32'h0;
memory[5395] <= 32'h0;
memory[5396] <= 32'h0;
memory[5397] <= 32'h0;
memory[5398] <= 32'h0;
memory[5399] <= 32'h0;
memory[5400] <= 32'h0;
memory[5401] <= 32'h0;
memory[5402] <= 32'h0;
memory[5403] <= 32'h0;
memory[5404] <= 32'h0;
memory[5405] <= 32'h0;
memory[5406] <= 32'h0;
memory[5407] <= 32'h0;
memory[5408] <= 32'h0;
memory[5409] <= 32'h0;
memory[5410] <= 32'h0;
memory[5411] <= 32'h0;
memory[5412] <= 32'h0;
memory[5413] <= 32'h0;
memory[5414] <= 32'h0;
memory[5415] <= 32'h0;
memory[5416] <= 32'h0;
memory[5417] <= 32'h0;
memory[5418] <= 32'h0;
memory[5419] <= 32'h0;
memory[5420] <= 32'h0;
memory[5421] <= 32'h0;
memory[5422] <= 32'h0;
memory[5423] <= 32'h0;
memory[5424] <= 32'h0;
memory[5425] <= 32'h0;
memory[5426] <= 32'h0;
memory[5427] <= 32'h0;
memory[5428] <= 32'h0;
memory[5429] <= 32'h0;
memory[5430] <= 32'h0;
memory[5431] <= 32'h0;
memory[5432] <= 32'h0;
memory[5433] <= 32'h0;
memory[5434] <= 32'h0;
memory[5435] <= 32'h0;
memory[5436] <= 32'h0;
memory[5437] <= 32'h0;
memory[5438] <= 32'h0;
memory[5439] <= 32'h0;
memory[5440] <= 32'h0;
memory[5441] <= 32'h0;
memory[5442] <= 32'h0;
memory[5443] <= 32'h0;
memory[5444] <= 32'h0;
memory[5445] <= 32'h0;
memory[5446] <= 32'h0;
memory[5447] <= 32'h0;
memory[5448] <= 32'h0;
memory[5449] <= 32'h0;
memory[5450] <= 32'h0;
memory[5451] <= 32'h0;
memory[5452] <= 32'h0;
memory[5453] <= 32'h0;
memory[5454] <= 32'h0;
memory[5455] <= 32'h0;
memory[5456] <= 32'h0;
memory[5457] <= 32'h0;
memory[5458] <= 32'h0;
memory[5459] <= 32'h0;
memory[5460] <= 32'h0;
memory[5461] <= 32'h0;
memory[5462] <= 32'h0;
memory[5463] <= 32'h0;
memory[5464] <= 32'h0;
memory[5465] <= 32'h0;
memory[5466] <= 32'h0;
memory[5467] <= 32'h0;
memory[5468] <= 32'h0;
memory[5469] <= 32'h0;
memory[5470] <= 32'h0;
memory[5471] <= 32'h0;
memory[5472] <= 32'h0;
memory[5473] <= 32'h0;
memory[5474] <= 32'h0;
memory[5475] <= 32'h0;
memory[5476] <= 32'h0;
memory[5477] <= 32'h0;
memory[5478] <= 32'h0;
memory[5479] <= 32'h0;
memory[5480] <= 32'h0;
memory[5481] <= 32'h0;
memory[5482] <= 32'h0;
memory[5483] <= 32'h0;
memory[5484] <= 32'h0;
memory[5485] <= 32'h0;
memory[5486] <= 32'h0;
memory[5487] <= 32'h0;
memory[5488] <= 32'h0;
memory[5489] <= 32'h0;
memory[5490] <= 32'h0;
memory[5491] <= 32'h0;
memory[5492] <= 32'h0;
memory[5493] <= 32'h0;
memory[5494] <= 32'h0;
memory[5495] <= 32'h0;
memory[5496] <= 32'h0;
memory[5497] <= 32'h0;
memory[5498] <= 32'h0;
memory[5499] <= 32'h0;
memory[5500] <= 32'h0;
memory[5501] <= 32'h0;
memory[5502] <= 32'h0;
memory[5503] <= 32'h0;
memory[5504] <= 32'h0;
memory[5505] <= 32'h0;
memory[5506] <= 32'h0;
memory[5507] <= 32'h0;
memory[5508] <= 32'h0;
memory[5509] <= 32'h0;
memory[5510] <= 32'h0;
memory[5511] <= 32'h0;
memory[5512] <= 32'h0;
memory[5513] <= 32'h0;
memory[5514] <= 32'h0;
memory[5515] <= 32'h0;
memory[5516] <= 32'h0;
memory[5517] <= 32'h0;
memory[5518] <= 32'h0;
memory[5519] <= 32'h0;
memory[5520] <= 32'h0;
memory[5521] <= 32'h0;
memory[5522] <= 32'h0;
memory[5523] <= 32'h0;
memory[5524] <= 32'h0;
memory[5525] <= 32'h0;
memory[5526] <= 32'h0;
memory[5527] <= 32'h0;
memory[5528] <= 32'h0;
memory[5529] <= 32'h0;
memory[5530] <= 32'h0;
memory[5531] <= 32'h0;
memory[5532] <= 32'h0;
memory[5533] <= 32'h0;
memory[5534] <= 32'h0;
memory[5535] <= 32'h0;
memory[5536] <= 32'h0;
memory[5537] <= 32'h0;
memory[5538] <= 32'h0;
memory[5539] <= 32'h0;
memory[5540] <= 32'h0;
memory[5541] <= 32'h0;
memory[5542] <= 32'h0;
memory[5543] <= 32'h0;
memory[5544] <= 32'h0;
memory[5545] <= 32'h0;
memory[5546] <= 32'h0;
memory[5547] <= 32'h0;
memory[5548] <= 32'h0;
memory[5549] <= 32'h0;
memory[5550] <= 32'h0;
memory[5551] <= 32'h0;
memory[5552] <= 32'h0;
memory[5553] <= 32'h0;
memory[5554] <= 32'h0;
memory[5555] <= 32'h0;
memory[5556] <= 32'h0;
memory[5557] <= 32'h0;
memory[5558] <= 32'h0;
memory[5559] <= 32'h0;
memory[5560] <= 32'h0;
memory[5561] <= 32'h0;
memory[5562] <= 32'h0;
memory[5563] <= 32'h0;
memory[5564] <= 32'h0;
memory[5565] <= 32'h0;
memory[5566] <= 32'h0;
memory[5567] <= 32'h0;
memory[5568] <= 32'h0;
memory[5569] <= 32'h0;
memory[5570] <= 32'h0;
memory[5571] <= 32'h0;
memory[5572] <= 32'h0;
memory[5573] <= 32'h0;
memory[5574] <= 32'h0;
memory[5575] <= 32'h0;
memory[5576] <= 32'h0;
memory[5577] <= 32'h0;
memory[5578] <= 32'h0;
memory[5579] <= 32'h0;
memory[5580] <= 32'h0;
memory[5581] <= 32'h0;
memory[5582] <= 32'h0;
memory[5583] <= 32'h0;
memory[5584] <= 32'h0;
memory[5585] <= 32'h0;
memory[5586] <= 32'h0;
memory[5587] <= 32'h0;
memory[5588] <= 32'h0;
memory[5589] <= 32'h0;
memory[5590] <= 32'h0;
memory[5591] <= 32'h0;
memory[5592] <= 32'h0;
memory[5593] <= 32'h0;
memory[5594] <= 32'h0;
memory[5595] <= 32'h0;
memory[5596] <= 32'h0;
memory[5597] <= 32'h0;
memory[5598] <= 32'h0;
memory[5599] <= 32'h0;
memory[5600] <= 32'h0;
memory[5601] <= 32'h0;
memory[5602] <= 32'h0;
memory[5603] <= 32'h0;
memory[5604] <= 32'h0;
memory[5605] <= 32'h0;
memory[5606] <= 32'h0;
memory[5607] <= 32'h0;
memory[5608] <= 32'h0;
memory[5609] <= 32'h0;
memory[5610] <= 32'h0;
memory[5611] <= 32'h0;
memory[5612] <= 32'h0;
memory[5613] <= 32'h0;
memory[5614] <= 32'h0;
memory[5615] <= 32'h0;
memory[5616] <= 32'h0;
memory[5617] <= 32'h0;
memory[5618] <= 32'h0;
memory[5619] <= 32'h0;
memory[5620] <= 32'h0;
memory[5621] <= 32'h0;
memory[5622] <= 32'h0;
memory[5623] <= 32'h0;
memory[5624] <= 32'h0;
memory[5625] <= 32'h0;
memory[5626] <= 32'h0;
memory[5627] <= 32'h0;
memory[5628] <= 32'h0;
memory[5629] <= 32'h0;
memory[5630] <= 32'h0;
memory[5631] <= 32'h0;
memory[5632] <= 32'h0;
memory[5633] <= 32'h0;
memory[5634] <= 32'h0;
memory[5635] <= 32'h0;
memory[5636] <= 32'h0;
memory[5637] <= 32'h0;
memory[5638] <= 32'h0;
memory[5639] <= 32'h0;
memory[5640] <= 32'h0;
memory[5641] <= 32'h0;
memory[5642] <= 32'h0;
memory[5643] <= 32'h0;
memory[5644] <= 32'h0;
memory[5645] <= 32'h0;
memory[5646] <= 32'h0;
memory[5647] <= 32'h0;
memory[5648] <= 32'h0;
memory[5649] <= 32'h0;
memory[5650] <= 32'h0;
memory[5651] <= 32'h0;
memory[5652] <= 32'h0;
memory[5653] <= 32'h0;
memory[5654] <= 32'h0;
memory[5655] <= 32'h0;
memory[5656] <= 32'h0;
memory[5657] <= 32'h0;
memory[5658] <= 32'h0;
memory[5659] <= 32'h0;
memory[5660] <= 32'h0;
memory[5661] <= 32'h0;
memory[5662] <= 32'h0;
memory[5663] <= 32'h0;
memory[5664] <= 32'h0;
memory[5665] <= 32'h0;
memory[5666] <= 32'h0;
memory[5667] <= 32'h0;
memory[5668] <= 32'h0;
memory[5669] <= 32'h0;
memory[5670] <= 32'h0;
memory[5671] <= 32'h0;
memory[5672] <= 32'h0;
memory[5673] <= 32'h0;
memory[5674] <= 32'h0;
memory[5675] <= 32'h0;
memory[5676] <= 32'h0;
memory[5677] <= 32'h0;
memory[5678] <= 32'h0;
memory[5679] <= 32'h0;
memory[5680] <= 32'h0;
memory[5681] <= 32'h0;
memory[5682] <= 32'h0;
memory[5683] <= 32'h0;
memory[5684] <= 32'h0;
memory[5685] <= 32'h0;
memory[5686] <= 32'h0;
memory[5687] <= 32'h0;
memory[5688] <= 32'h0;
memory[5689] <= 32'h0;
memory[5690] <= 32'h0;
memory[5691] <= 32'h0;
memory[5692] <= 32'h0;
memory[5693] <= 32'h0;
memory[5694] <= 32'h0;
memory[5695] <= 32'h0;
memory[5696] <= 32'h0;
memory[5697] <= 32'h0;
memory[5698] <= 32'h0;
memory[5699] <= 32'h0;
memory[5700] <= 32'h0;
memory[5701] <= 32'h0;
memory[5702] <= 32'h0;
memory[5703] <= 32'h0;
memory[5704] <= 32'h0;
memory[5705] <= 32'h0;
memory[5706] <= 32'h0;
memory[5707] <= 32'h0;
memory[5708] <= 32'h0;
memory[5709] <= 32'h0;
memory[5710] <= 32'h0;
memory[5711] <= 32'h0;
memory[5712] <= 32'h0;
memory[5713] <= 32'h0;
memory[5714] <= 32'h0;
memory[5715] <= 32'h0;
memory[5716] <= 32'h0;
memory[5717] <= 32'h0;
memory[5718] <= 32'h0;
memory[5719] <= 32'h0;
memory[5720] <= 32'h0;
memory[5721] <= 32'h0;
memory[5722] <= 32'h0;
memory[5723] <= 32'h0;
memory[5724] <= 32'h0;
memory[5725] <= 32'h0;
memory[5726] <= 32'h0;
memory[5727] <= 32'h0;
memory[5728] <= 32'h0;
memory[5729] <= 32'h0;
memory[5730] <= 32'h0;
memory[5731] <= 32'h0;
memory[5732] <= 32'h0;
memory[5733] <= 32'h0;
memory[5734] <= 32'h0;
memory[5735] <= 32'h0;
memory[5736] <= 32'h0;
memory[5737] <= 32'h0;
memory[5738] <= 32'h0;
memory[5739] <= 32'h0;
memory[5740] <= 32'h0;
memory[5741] <= 32'h0;
memory[5742] <= 32'h0;
memory[5743] <= 32'h0;
memory[5744] <= 32'h0;
memory[5745] <= 32'h0;
memory[5746] <= 32'h0;
memory[5747] <= 32'h0;
memory[5748] <= 32'h0;
memory[5749] <= 32'h0;
memory[5750] <= 32'h0;
memory[5751] <= 32'h0;
memory[5752] <= 32'h0;
memory[5753] <= 32'h0;
memory[5754] <= 32'h0;
memory[5755] <= 32'h0;
memory[5756] <= 32'h0;
memory[5757] <= 32'h0;
memory[5758] <= 32'h0;
memory[5759] <= 32'h0;
memory[5760] <= 32'h0;
memory[5761] <= 32'h0;
memory[5762] <= 32'h0;
memory[5763] <= 32'h0;
memory[5764] <= 32'h0;
memory[5765] <= 32'h0;
memory[5766] <= 32'h0;
memory[5767] <= 32'h0;
memory[5768] <= 32'h0;
memory[5769] <= 32'h0;
memory[5770] <= 32'h0;
memory[5771] <= 32'h0;
memory[5772] <= 32'h0;
memory[5773] <= 32'h0;
memory[5774] <= 32'h0;
memory[5775] <= 32'h0;
memory[5776] <= 32'h0;
memory[5777] <= 32'h0;
memory[5778] <= 32'h0;
memory[5779] <= 32'h0;
memory[5780] <= 32'h0;
memory[5781] <= 32'h0;
memory[5782] <= 32'h0;
memory[5783] <= 32'h0;
memory[5784] <= 32'h0;
memory[5785] <= 32'h0;
memory[5786] <= 32'h0;
memory[5787] <= 32'h0;
memory[5788] <= 32'h0;
memory[5789] <= 32'h0;
memory[5790] <= 32'h0;
memory[5791] <= 32'h0;
memory[5792] <= 32'h0;
memory[5793] <= 32'h0;
memory[5794] <= 32'h0;
memory[5795] <= 32'h0;
memory[5796] <= 32'h0;
memory[5797] <= 32'h0;
memory[5798] <= 32'h0;
memory[5799] <= 32'h0;
memory[5800] <= 32'h0;
memory[5801] <= 32'h0;
memory[5802] <= 32'h0;
memory[5803] <= 32'h0;
memory[5804] <= 32'h0;
memory[5805] <= 32'h0;
memory[5806] <= 32'h0;
memory[5807] <= 32'h0;
memory[5808] <= 32'h0;
memory[5809] <= 32'h0;
memory[5810] <= 32'h0;
memory[5811] <= 32'h0;
memory[5812] <= 32'h0;
memory[5813] <= 32'h0;
memory[5814] <= 32'h0;
memory[5815] <= 32'h0;
memory[5816] <= 32'h0;
memory[5817] <= 32'h0;
memory[5818] <= 32'h0;
memory[5819] <= 32'h0;
memory[5820] <= 32'h0;
memory[5821] <= 32'h0;
memory[5822] <= 32'h0;
memory[5823] <= 32'h0;
memory[5824] <= 32'h0;
memory[5825] <= 32'h0;
memory[5826] <= 32'h0;
memory[5827] <= 32'h0;
memory[5828] <= 32'h0;
memory[5829] <= 32'h0;
memory[5830] <= 32'h0;
memory[5831] <= 32'h0;
memory[5832] <= 32'h0;
memory[5833] <= 32'h0;
memory[5834] <= 32'h0;
memory[5835] <= 32'h0;
memory[5836] <= 32'h0;
memory[5837] <= 32'h0;
memory[5838] <= 32'h0;
memory[5839] <= 32'h0;
memory[5840] <= 32'h0;
memory[5841] <= 32'h0;
memory[5842] <= 32'h0;
memory[5843] <= 32'h0;
memory[5844] <= 32'h0;
memory[5845] <= 32'h0;
memory[5846] <= 32'h0;
memory[5847] <= 32'h0;
memory[5848] <= 32'h0;
memory[5849] <= 32'h0;
memory[5850] <= 32'h0;
memory[5851] <= 32'h0;
memory[5852] <= 32'h0;
memory[5853] <= 32'h0;
memory[5854] <= 32'h0;
memory[5855] <= 32'h0;
memory[5856] <= 32'h0;
memory[5857] <= 32'h0;
memory[5858] <= 32'h0;
memory[5859] <= 32'h0;
memory[5860] <= 32'h0;
memory[5861] <= 32'h0;
memory[5862] <= 32'h0;
memory[5863] <= 32'h0;
memory[5864] <= 32'h0;
memory[5865] <= 32'h0;
memory[5866] <= 32'h0;
memory[5867] <= 32'h0;
memory[5868] <= 32'h0;
memory[5869] <= 32'h0;
memory[5870] <= 32'h0;
memory[5871] <= 32'h0;
memory[5872] <= 32'h0;
memory[5873] <= 32'h0;
memory[5874] <= 32'h0;
memory[5875] <= 32'h0;
memory[5876] <= 32'h0;
memory[5877] <= 32'h0;
memory[5878] <= 32'h0;
memory[5879] <= 32'h1;
memory[5880] <= 32'h1;
memory[5881] <= 32'h1;
memory[5882] <= 32'h1;
memory[5883] <= 32'h0;
memory[5884] <= 32'h0;
memory[5885] <= 32'h0;
memory[5886] <= 32'h0;
memory[5887] <= 32'h0;
memory[5888] <= 32'h0;
memory[5889] <= 32'h0;
memory[5890] <= 32'h0;
memory[5891] <= 32'h0;
memory[5892] <= 32'h0;
memory[5893] <= 32'h0;
memory[5894] <= 32'h0;
memory[5895] <= 32'h0;
memory[5896] <= 32'h0;
memory[5897] <= 32'h0;
memory[5898] <= 32'h0;
memory[5899] <= 32'h0;
memory[5900] <= 32'h0;
memory[5901] <= 32'h0;
memory[5902] <= 32'h0;
memory[5903] <= 32'h0;
memory[5904] <= 32'h0;
memory[5905] <= 32'h0;
memory[5906] <= 32'h0;
memory[5907] <= 32'h0;
memory[5908] <= 32'h0;
memory[5909] <= 32'h0;
memory[5910] <= 32'h0;
memory[5911] <= 32'h1;
memory[5912] <= 32'h1;
memory[5913] <= 32'h1;
memory[5914] <= 32'h1;
memory[5915] <= 32'h0;
memory[5916] <= 32'h0;
memory[5917] <= 32'h0;
memory[5918] <= 32'h0;
memory[5919] <= 32'h0;
memory[5920] <= 32'h0;
memory[5921] <= 32'h0;
memory[5922] <= 32'h0;
memory[5923] <= 32'h0;
memory[5924] <= 32'h0;
memory[5925] <= 32'h0;
memory[5926] <= 32'h0;
memory[5927] <= 32'h0;
memory[5928] <= 32'h0;
memory[5929] <= 32'h0;
memory[5930] <= 32'h0;
memory[5931] <= 32'h0;
memory[5932] <= 32'h0;
memory[5933] <= 32'h0;
memory[5934] <= 32'h0;
memory[5935] <= 32'h0;
memory[5936] <= 32'h0;
memory[5937] <= 32'h0;
memory[5938] <= 32'h0;
memory[5939] <= 32'h0;
memory[5940] <= 32'h0;
memory[5941] <= 32'h0;
memory[5942] <= 32'h0;
memory[5943] <= 32'h1;
memory[5944] <= 32'h1;
memory[5945] <= 32'h1;
memory[5946] <= 32'h1;
memory[5947] <= 32'h0;
memory[5948] <= 32'h0;
memory[5949] <= 32'h0;
memory[5950] <= 32'h0;
memory[5951] <= 32'h0;
memory[5952] <= 32'h0;
memory[5953] <= 32'h0;
memory[5954] <= 32'h0;
memory[5955] <= 32'h0;
memory[5956] <= 32'h0;
memory[5957] <= 32'h0;
memory[5958] <= 32'h0;
memory[5959] <= 32'h0;
memory[5960] <= 32'h0;
memory[5961] <= 32'h0;
memory[5962] <= 32'h0;
memory[5963] <= 32'h0;
memory[5964] <= 32'h0;
memory[5965] <= 32'h0;
memory[5966] <= 32'h0;
memory[5967] <= 32'h0;
memory[5968] <= 32'h0;
memory[5969] <= 32'h0;
memory[5970] <= 32'h0;
memory[5971] <= 32'h0;
memory[5972] <= 32'h0;
memory[5973] <= 32'h0;
memory[5974] <= 32'h0;
memory[5975] <= 32'h1;
memory[5976] <= 32'h1;
memory[5977] <= 32'h1;
memory[5978] <= 32'h1;
memory[5979] <= 32'h0;
memory[5980] <= 32'h0;
memory[5981] <= 32'h0;
memory[5982] <= 32'h0;
memory[5983] <= 32'h0;
memory[5984] <= 32'h0;
memory[5985] <= 32'h0;
memory[5986] <= 32'h0;
memory[5987] <= 32'h0;
memory[5988] <= 32'h0;
memory[5989] <= 32'h0;
memory[5990] <= 32'h0;
memory[5991] <= 32'h0;
memory[5992] <= 32'h0;
memory[5993] <= 32'h0;
memory[5994] <= 32'h0;
memory[5995] <= 32'h0;
memory[5996] <= 32'h0;
memory[5997] <= 32'h0;
memory[5998] <= 32'h0;
memory[5999] <= 32'h0;
memory[6000] <= 32'h0;
memory[6001] <= 32'h0;
memory[6002] <= 32'h0;
memory[6003] <= 32'h0;
memory[6004] <= 32'h0;
memory[6005] <= 32'h0;
memory[6006] <= 32'h0;
memory[6007] <= 32'h1;
memory[6008] <= 32'h1;
memory[6009] <= 32'h1;
memory[6010] <= 32'h1;
memory[6011] <= 32'h0;
memory[6012] <= 32'h0;
memory[6013] <= 32'h0;
memory[6014] <= 32'h0;
memory[6015] <= 32'h0;
memory[6016] <= 32'h0;
memory[6017] <= 32'h0;
memory[6018] <= 32'h0;
memory[6019] <= 32'h0;
memory[6020] <= 32'h0;
memory[6021] <= 32'h0;
memory[6022] <= 32'h0;
memory[6023] <= 32'h0;
memory[6024] <= 32'h0;
memory[6025] <= 32'h0;
memory[6026] <= 32'h0;
memory[6027] <= 32'h0;
memory[6028] <= 32'h0;
memory[6029] <= 32'h0;
memory[6030] <= 32'h0;
memory[6031] <= 32'h0;
memory[6032] <= 32'h0;
memory[6033] <= 32'h0;
memory[6034] <= 32'h0;
memory[6035] <= 32'h0;
memory[6036] <= 32'h0;
memory[6037] <= 32'h0;
memory[6038] <= 32'h0;
memory[6039] <= 32'h1;
memory[6040] <= 32'h1;
memory[6041] <= 32'h1;
memory[6042] <= 32'h1;
memory[6043] <= 32'h0;
memory[6044] <= 32'h0;
memory[6045] <= 32'h0;
memory[6046] <= 32'h0;
memory[6047] <= 32'h0;
memory[6048] <= 32'h0;
memory[6049] <= 32'h0;
memory[6050] <= 32'h0;
memory[6051] <= 32'h0;
memory[6052] <= 32'h0;
memory[6053] <= 32'h0;
memory[6054] <= 32'h0;
memory[6055] <= 32'h0;
memory[6056] <= 32'h0;
memory[6057] <= 32'h0;
memory[6058] <= 32'h0;
memory[6059] <= 32'h0;
memory[6060] <= 32'h0;
memory[6061] <= 32'h0;
memory[6062] <= 32'h0;
memory[6063] <= 32'h0;
memory[6064] <= 32'h0;
memory[6065] <= 32'h0;
memory[6066] <= 32'h0;
memory[6067] <= 32'h0;
memory[6068] <= 32'h0;
memory[6069] <= 32'h0;
memory[6070] <= 32'h0;
memory[6071] <= 32'h1;
memory[6072] <= 32'h1;
memory[6073] <= 32'h1;
memory[6074] <= 32'h1;
memory[6075] <= 32'h0;
memory[6076] <= 32'h0;
memory[6077] <= 32'h0;
memory[6078] <= 32'h0;
memory[6079] <= 32'h0;
memory[6080] <= 32'h0;
memory[6081] <= 32'h0;
memory[6082] <= 32'h0;
memory[6083] <= 32'h0;
memory[6084] <= 32'h0;
memory[6085] <= 32'h0;
memory[6086] <= 32'h0;
memory[6087] <= 32'h0;
memory[6088] <= 32'h0;
memory[6089] <= 32'h0;
memory[6090] <= 32'h0;
memory[6091] <= 32'h0;
memory[6092] <= 32'h0;
memory[6093] <= 32'h0;
memory[6094] <= 32'h0;
memory[6095] <= 32'h0;
memory[6096] <= 32'h0;
memory[6097] <= 32'h0;
memory[6098] <= 32'h0;
memory[6099] <= 32'h0;
memory[6100] <= 32'h0;
memory[6101] <= 32'h0;
memory[6102] <= 32'h0;
memory[6103] <= 32'h1;
memory[6104] <= 32'h1;
memory[6105] <= 32'h1;
memory[6106] <= 32'h1;
memory[6107] <= 32'h1;
memory[6108] <= 32'h1;
memory[6109] <= 32'h1;
memory[6110] <= 32'h1;
memory[6111] <= 32'h1;
memory[6112] <= 32'h1;
memory[6113] <= 32'h1;
memory[6114] <= 32'h1;
memory[6115] <= 32'h1;
memory[6116] <= 32'h1;
memory[6117] <= 32'h1;
memory[6118] <= 32'h1;
memory[6119] <= 32'h1;
memory[6120] <= 32'h1;
memory[6121] <= 32'h1;
memory[6122] <= 32'h1;
memory[6123] <= 32'h1;
memory[6124] <= 32'h1;
memory[6125] <= 32'h1;
memory[6126] <= 32'h1;
memory[6127] <= 32'h1;
memory[6128] <= 32'h1;
memory[6129] <= 32'h1;
memory[6130] <= 32'h1;
memory[6131] <= 32'h1;
memory[6132] <= 32'h1;
memory[6133] <= 32'h1;
memory[6134] <= 32'h1;
memory[6135] <= 32'h1;
memory[6136] <= 32'h1;
memory[6137] <= 32'h1;
memory[6138] <= 32'h1;
memory[6139] <= 32'h0;





 
    end
   
    always @(posedge Clk) 
    begin
        if (MemWrite)   
        begin                           
            if(whb == 2'b0)
            begin
                memory[Address[15:2]] <= WriteData;
            end
            
            else if(whb == 2'b01)
            begin
                memory[Address[15:2]] <= {16'b0,WriteData[15:0]};
            end
                
            else if(whb == 2'b10)
            begin
                memory[Address[15:2]] <= {24'b0,WriteData[7:0]};
            end
        end
    end
    
    always @(*) 
    begin
        if (MemRead)   
        begin                           
            if(whb == 2'b0)
            begin
                ReadData <= memory[Address[15:2]];
            end
            
            else if(whb == 2'b01)
            begin
                if(memory[Address[15:2]][15] == 0) begin
                    ReadData <= {16'b0,memory[Address[15:2]][15:0]};
                end
                else begin
                    ReadData <= {16'b1111111111111111,memory[Address[15:2]][15:0]};
                end
            end
                
            else if(whb == 2'b10)
            begin
                if(memory[Address[11:2]][7] == 0) begin
                    ReadData <= {24'b0,memory[Address[15:2]][7:0]};
                end
                else begin
                    ReadData <= {24'b111111111111111111111111,memory[Address[15:2]][7:0]};
                end
            end
        end
    end
endmodule
